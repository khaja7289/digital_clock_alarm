* NGSPICE file created from alarm_clock_top.ext - technology: scmos

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 Q CLK D gnd vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

.subckt alarm_clock_top vdd gnd clock key[0] key[1] key[2] key[3] reset time_button
+ alarm_button fastwatch ms_hour[0] ms_hour[1] ms_hour[2] ms_hour[3] ms_hour[4] ms_hour[5]
+ ms_hour[6] ms_hour[7] ls_hour[0] ls_hour[1] ls_hour[2] ls_hour[3] ls_hour[4] ls_hour[5]
+ ls_hour[6] ls_hour[7] ms_minute[0] ms_minute[1] ms_minute[2] ms_minute[3] ms_minute[4]
+ ms_minute[5] ms_minute[6] ms_minute[7] ls_minute[0] ls_minute[1] ls_minute[2] ls_minute[3]
+ ls_minute[4] ls_minute[5] ls_minute[6] ls_minute[7] alarm_sound
XAND2X2_5 INVX1_31/Y AND2X2_5/B gnd AND2X2_5/Y vdd AND2X2
XMUX2X1_17 MUX2X1_33/A MUX2X1_5/A AND2X2_4/Y gnd NOR2X1_69/B vdd MUX2X1
XMUX2X1_39 MUX2X1_2/A MUX2X1_39/B BUFX4_4/Y gnd MUX2X1_39/Y vdd MUX2X1
XMUX2X1_28 MUX2X1_46/A MUX2X1_34/A AND2X2_4/Y gnd NOR2X1_80/B vdd MUX2X1
XNAND2X1_43 MUX2X1_6/B BUFX4_9/Y gnd OAI21X1_57/C vdd NAND2X1
XNAND2X1_32 NOR3X1_9/Y NOR3X1_11/Y gnd NOR2X1_85/A vdd NAND2X1
XNAND2X1_54 NAND3X1_1/B OAI21X1_2/A gnd OR2X2_1/A vdd NAND2X1
XNAND2X1_21 INVX2_8/A NOR3X1_7/B gnd NOR3X1_8/C vdd NAND2X1
XNAND2X1_10 XOR2X1_8/B NOR2X1_32/Y gnd NAND3X1_4/C vdd NAND2X1
XOAI22X1_3 OAI22X1_3/A OAI22X1_3/B OAI22X1_3/C OAI22X1_3/D gnd OAI22X1_3/Y vdd OAI22X1
XINVX2_12 INVX2_12/A gnd INVX2_12/Y vdd INVX2
XOAI21X1_19 INVX1_11/Y INVX2_4/Y BUFX4_13/Y gnd OAI21X1_19/Y vdd OAI21X1
XFILL_11_1_0 gnd vdd FILL
XFILL_3_2_0 gnd vdd FILL
XDFFPOSX1_125 MUX2X1_3/A NOR2X1_75/A NOR2X1_75/Y gnd vdd DFFPOSX1
XDFFPOSX1_136 MUX2X1_35/A CLKBUF1_1/Y NOR2X1_78/Y gnd vdd DFFPOSX1
XDFFPOSX1_103 INVX2_12/A CLKBUF1_2/Y NOR2X1_54/Y gnd vdd DFFPOSX1
XDFFPOSX1_114 INVX2_8/A NOR2X1_104/A AOI21X1_31/Y gnd vdd DFFPOSX1
XDFFPOSX1_147 MUX2X1_9/A CLKBUF1_5/Y NOR2X1_81/Y gnd vdd DFFPOSX1
XXNOR2X1_6 XNOR2X1_6/A INVX2_12/Y gnd XNOR2X1_6/Y vdd XNOR2X1
XFILL_0_0_0 gnd vdd FILL
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XOR2X2_4 OR2X2_4/A time_button gnd OR2X2_4/Y vdd OR2X2
XFILL_16_0_0 gnd vdd FILL
XFILL_8_1_0 gnd vdd FILL
XAND2X2_6 INVX2_14/Y AND2X2_6/B gnd AND2X2_6/Y vdd AND2X2
XMUX2X1_18 MUX2X1_35/A MUX2X1_6/A AND2X2_4/Y gnd NOR2X1_70/B vdd MUX2X1
XMUX2X1_29 MUX2X1_1/A MUX2X1_9/A AND2X2_4/Y gnd NOR2X1_81/B vdd MUX2X1
XNAND2X1_11 INVX2_4/A INVX1_11/Y gnd OR2X2_3/A vdd NAND2X1
XNAND2X1_44 XOR2X1_6/A BUFX4_8/Y gnd OAI21X1_58/C vdd NAND2X1
XNAND2X1_55 INVX2_10/A fastwatch gnd OAI21X1_66/C vdd NAND2X1
XNAND2X1_33 NOR3X1_12/Y NOR3X1_10/Y gnd NOR2X1_85/B vdd NAND2X1
XAOI22X1_1 AOI22X1_1/A NOR3X1_7/Y NOR3X1_5/Y AOI22X1_1/D gnd AOI22X1_1/Y vdd AOI22X1
XNAND2X1_22 INVX2_8/Y NOR3X1_5/C gnd NOR2X1_47/B vdd NAND2X1
XOAI22X1_4 OAI22X1_4/A OAI22X1_4/B OAI22X1_4/C OAI22X1_4/D gnd OAI22X1_4/Y vdd OAI22X1
XFILL_11_1_1 gnd vdd FILL
XFILL_3_2_1 gnd vdd FILL
XINVX2_13 INVX2_13/A gnd INVX2_13/Y vdd INVX2
XDFFPOSX1_126 MUX2X1_4/A NOR2X1_77/A NOR2X1_76/Y gnd vdd DFFPOSX1
XDFFPOSX1_137 MUX2X1_36/A CLKBUF1_1/Y NOR2X1_79/Y gnd vdd DFFPOSX1
XDFFPOSX1_148 MUX2X1_47/A CLKBUF1_5/Y NOR2X1_82/Y gnd vdd DFFPOSX1
XDFFPOSX1_104 INVX1_22/A CLKBUF1_2/Y AOI21X1_26/Y gnd vdd DFFPOSX1
XDFFPOSX1_115 INVX2_9/A NOR2X1_23/A AOI21X1_32/Y gnd vdd DFFPOSX1
XFILL_10_1 gnd vdd FILL
XFILL_0_0_1 gnd vdd FILL
XOR2X2_5 time_button OR2X2_5/B gnd OR2X2_5/Y vdd OR2X2
XXNOR2X1_7 XNOR2X1_7/A INVX2_13/Y gnd XNOR2X1_7/Y vdd XNOR2X1
XFILL_16_0_1 gnd vdd FILL
XFILL_8_1_1 gnd vdd FILL
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XAND2X2_7 INVX2_14/Y AND2X2_7/B gnd AND2X2_7/Y vdd AND2X2
XMUX2X1_19 MUX2X1_36/A MUX2X1_7/A AND2X2_4/Y gnd NOR2X1_71/B vdd MUX2X1
XNAND2X1_12 OAI21X1_21/Y OR2X2_3/Y gnd NAND2X1_12/Y vdd NAND2X1
XNAND2X1_34 NOR2X1_86/A BUFX4_5/Y gnd OAI21X1_46/C vdd NAND2X1
XNAND2X1_45 XOR2X1_5/A BUFX4_9/Y gnd OAI21X1_59/C vdd NAND2X1
XNAND2X1_56 AND2X2_19/Y AOI21X1_4/A gnd OAI21X1_5/B vdd NAND2X1
XNAND2X1_23 NOR3X1_7/B INVX2_8/Y gnd NOR2X1_48/B vdd NAND2X1
XAOI22X1_2 AOI22X1_2/A NOR3X1_7/Y OR2X2_9/Y AND2X2_4/A gnd AOI22X1_2/Y vdd AOI22X1
XINVX2_14 alarm_button gnd INVX2_14/Y vdd INVX2
XDFFPOSX1_127 MUX2X1_5/A NOR2X1_77/A NOR2X1_69/Y gnd vdd DFFPOSX1
XDFFPOSX1_116 NOR3X1_7/B CLKBUF1_6/Y AOI21X1_29/Y gnd vdd DFFPOSX1
XDFFPOSX1_105 INVX1_23/A INVX2_11/A NOR2X1_59/Y gnd vdd DFFPOSX1
XDFFPOSX1_138 MUX2X1_34/A CLKBUF1_5/Y NOR2X1_80/Y gnd vdd DFFPOSX1
XDFFPOSX1_149 MUX2X1_48/A CLKBUF1_5/Y NOR2X1_83/Y gnd vdd DFFPOSX1
XBUFX4_10 INVX8_1/Y gnd BUFX4_10/Y vdd BUFX4
XINVX8_1 INVX8_1/A gnd INVX8_1/Y vdd INVX8
XOR2X2_6 alarm_button OR2X2_6/B gnd OR2X2_6/Y vdd OR2X2
XINVX1_8 INVX1_8/A gnd OR2X2_3/B vdd INVX1
XFILL_9_1 gnd vdd FILL
XAND2X2_8 INVX1_26/A BUFX2_56/A gnd BUFX2_50/A vdd AND2X2
XAOI22X1_3 BUFX4_6/Y AOI22X1_3/B NOR3X1_5/Y AOI22X1_3/D gnd AOI22X1_3/Y vdd AOI22X1
XNAND2X1_13 INVX4_1/A INVX1_12/Y gnd NOR3X1_3/A vdd NAND2X1
XNAND2X1_35 NOR2X1_87/A BUFX4_8/Y gnd OAI21X1_47/C vdd NAND2X1
XNAND2X1_57 INVX1_3/A INVX1_2/A gnd INVX1_4/A vdd NAND2X1
XNOR3X1_1 NOR3X1_1/A NOR3X1_1/B NOR3X1_1/C gnd NOR3X1_1/Y vdd NOR3X1
XNAND2X1_46 MUX2X1_9/B BUFX4_7/Y gnd OAI21X1_61/C vdd NAND2X1
XNAND2X1_24 INVX2_11/Y NOR3X1_6/Y gnd NOR2X1_54/B vdd NAND2X1
XFILL_6_2_0 gnd vdd FILL
XFILL_14_1_0 gnd vdd FILL
XINVX2_15 INVX2_15/A gnd INVX2_15/Y vdd INVX2
XDFFPOSX1_139 MUX2X1_1/A CLKBUF1_2/Y NOR2X1_73/Y gnd vdd DFFPOSX1
XDFFPOSX1_128 MUX2X1_6/A NOR2X1_79/A NOR2X1_70/Y gnd vdd DFFPOSX1
XDFFPOSX1_117 INVX2_8/A CLKBUF1_6/Y AOI21X1_31/Y gnd vdd DFFPOSX1
XDFFPOSX1_106 INVX1_24/A NOR2X1_104/A NOR2X1_60/Y gnd vdd DFFPOSX1
XFILL_3_0_0 gnd vdd FILL
XINVX8_2 INVX8_2/A gnd INVX8_2/Y vdd INVX8
XBUFX4_11 INVX8_1/Y gnd BUFX4_11/Y vdd BUFX4
XOR2X2_7 OR2X2_7/A OR2X2_7/B gnd OR2X2_7/Y vdd OR2X2
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XFILL_9_2 gnd vdd FILL
XAND2X2_9 NOR3X1_7/Y INVX2_14/Y gnd AND2X2_9/Y vdd AND2X2
XAOI22X1_4 AOI22X1_4/A NOR3X1_7/Y OR2X2_9/Y AND2X2_4/A gnd AOI22X1_4/Y vdd AOI22X1
XNAND2X1_14 XOR2X1_1/B INVX2_5/Y gnd NOR3X1_3/C vdd NAND2X1
XNAND2X1_36 XOR2X1_2/A BUFX4_8/Y gnd OAI21X1_48/C vdd NAND2X1
XNAND2X1_25 XNOR2X1_6/A OAI21X1_41/Y gnd NOR2X1_53/A vdd NAND2X1
XNAND2X1_58 INVX1_6/A AOI21X1_8/C gnd NOR3X1_2/B vdd NAND2X1
XNOR3X1_2 NOR3X1_2/A NOR3X1_2/B NOR3X1_2/C gnd NOR3X1_2/Y vdd NOR3X1
XNAND2X1_47 NOR2X1_99/A BUFX4_7/Y gnd OAI21X1_62/C vdd NAND2X1
XFILL_14_1_1 gnd vdd FILL
XFILL_6_2_1 gnd vdd FILL
XINVX2_16 NOR2X1_6/A gnd NOR3X1_2/A vdd INVX2
XDFFPOSX1_129 MUX2X1_7/A NOR2X1_79/A NOR2X1_71/Y gnd vdd DFFPOSX1
XCLKBUF1_1 clock gnd CLKBUF1_1/Y vdd CLKBUF1
XDFFPOSX1_118 INVX2_9/A CLKBUF1_6/Y AOI21X1_32/Y gnd vdd DFFPOSX1
XDFFPOSX1_107 INVX2_13/A NOR2X1_104/A NOR2X1_61/Y gnd vdd DFFPOSX1
XFILL_3_0_1 gnd vdd FILL
XBUFX4_12 INVX8_1/Y gnd BUFX4_12/Y vdd BUFX4
XOR2X2_8 alarm_button OR2X2_8/B gnd OR2X2_8/Y vdd OR2X2
XNAND2X1_15 INVX2_5/Y INVX1_13/Y gnd NOR2X1_38/A vdd NAND2X1
XNAND2X1_37 XOR2X1_1/A BUFX4_6/Y gnd OAI21X1_49/C vdd NAND2X1
XNAND2X1_26 INVX1_22/Y NOR2X1_55/Y gnd NAND2X1_26/Y vdd NAND2X1
XNAND2X1_59 AND2X2_2/B NOR3X1_2/A gnd NOR2X1_106/B vdd NAND2X1
XNAND2X1_48 XOR2X1_8/A BUFX4_7/Y gnd OAI21X1_63/C vdd NAND2X1
XNOR3X1_3 NOR3X1_3/A NOR3X1_3/B NOR3X1_3/C gnd NOR3X1_3/Y vdd NOR3X1
XINVX2_17 OR2X2_10/A gnd INVX2_17/Y vdd INVX2
XDFFPOSX1_119 MUX2X1_33/A NOR2X1_77/A NOR2X1_77/Y gnd vdd DFFPOSX1
XCLKBUF1_2 clock gnd CLKBUF1_2/Y vdd CLKBUF1
XMUX2X1_1 MUX2X1_1/A MUX2X1_1/B MUX2X1_9/S gnd MUX2X1_1/Y vdd MUX2X1
XDFFPOSX1_108 INVX1_25/A INVX8_2/A AOI21X1_27/Y gnd vdd DFFPOSX1
XBUFX4_13 INVX8_1/Y gnd BUFX4_13/Y vdd BUFX4
XDFFPOSX1_90 INVX1_48/A CLKBUF1_3/Y AOI21X1_23/Y gnd vdd DFFPOSX1
XOR2X2_9 OR2X2_9/A OR2X2_9/B gnd OR2X2_9/Y vdd OR2X2
XFILL_12_2_0 gnd vdd FILL
XFILL_7_1 gnd vdd FILL
XFILL_1_1_0 gnd vdd FILL
XNAND3X1_1 INVX1_4/Y NAND3X1_1/B OAI21X1_2/A gnd NOR3X1_2/C vdd NAND3X1
XNAND2X1_16 INVX2_5/A NOR2X1_35/Y gnd INVX1_14/A vdd NAND2X1
XNAND2X1_38 MUX2X1_1/B BUFX4_5/Y gnd OAI21X1_51/C vdd NAND2X1
XFILL_9_2_0 gnd vdd FILL
XNAND2X1_27 INVX2_11/Y NOR3X1_5/Y gnd NOR2X1_61/A vdd NAND2X1
XNAND2X1_49 XOR2X1_7/A BUFX4_6/Y gnd OAI21X1_64/C vdd NAND2X1
XNOR3X1_4 OR2X2_2/A NOR3X1_4/B NOR3X1_4/C gnd NOR3X1_4/Y vdd NOR3X1
XMUX2X1_2 MUX2X1_2/A MUX2X1_2/B MUX2X1_9/S gnd MUX2X1_2/Y vdd MUX2X1
XCLKBUF1_3 clock gnd CLKBUF1_3/Y vdd CLKBUF1
XXOR2X1_1 XOR2X1_1/A XOR2X1_1/B gnd XOR2X1_1/Y vdd XOR2X1
XDFFPOSX1_109 INVX1_23/A CLKBUF1_4/Y NOR2X1_59/Y gnd vdd DFFPOSX1
XFILL_6_0_0 gnd vdd FILL
XDFFPOSX1_91 INVX2_7/A CLKBUF1_3/Y AOI21X1_24/Y gnd vdd DFFPOSX1
XDFFPOSX1_80 INVX1_9/A NOR2X1_23/A NOR2X1_33/Y gnd vdd DFFPOSX1
XBUFX4_14 INVX8_1/Y gnd BUFX4_14/Y vdd BUFX4
XFILL_12_2_1 gnd vdd FILL
XFILL_7_2 gnd vdd FILL
XNAND3X1_2 INVX1_41/A XNOR2X1_2/B INVX2_4/Y gnd NOR2X1_30/B vdd NAND3X1
XNAND2X1_39 MUX2X1_2/B BUFX4_5/Y gnd OAI21X1_52/C vdd NAND2X1
XFILL_9_2_1 gnd vdd FILL
XNAND2X1_17 NOR2X1_39/Y NOR2X1_40/Y gnd NOR3X1_4/B vdd NAND2X1
XFILL_1_1_1 gnd vdd FILL
XNAND2X1_28 XNOR2X1_7/A OAI21X1_44/Y gnd NOR2X1_60/A vdd NAND2X1
XNOR3X1_5 INVX2_8/A INVX2_9/A NOR3X1_5/C gnd NOR3X1_5/Y vdd NOR3X1
XMUX2X1_3 MUX2X1_3/A XOR2X1_4/A MUX2X1_9/S gnd MUX2X1_3/Y vdd MUX2X1
XXOR2X1_2 XOR2X1_2/A INVX2_5/A gnd XOR2X1_2/Y vdd XOR2X1
XCLKBUF1_4 clock gnd CLKBUF1_4/Y vdd CLKBUF1
XFILL_6_0_1 gnd vdd FILL
XDFFPOSX1_81 INVX4_1/A CLKBUF1_1/Y AOI21X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_70 INVX2_4/A NOR2X1_75/A NOR2X1_34/Y gnd vdd DFFPOSX1
XDFFPOSX1_92 XOR2X1_5/B CLKBUF1_8/Y AOI21X1_25/Y gnd vdd DFFPOSX1
XNAND3X1_3 NAND3X1_3/A XNOR2X1_3/A OR2X2_2/Y gnd NAND3X1_3/Y vdd NAND3X1
XNAND2X1_18 INVX2_6/A INVX1_48/A gnd NOR3X1_3/B vdd NAND2X1
XNOR3X1_6 INVX2_8/Y NOR3X1_7/B OR2X2_9/A gnd NOR3X1_6/Y vdd NOR3X1
XNAND2X1_29 INVX1_25/Y NOR2X1_62/Y gnd NAND2X1_29/Y vdd NAND2X1
XMUX2X1_4 MUX2X1_4/A XOR2X1_3/A MUX2X1_9/S gnd MUX2X1_4/Y vdd MUX2X1
XXOR2X1_3 XOR2X1_3/A INVX2_3/A gnd XOR2X1_3/Y vdd XOR2X1
XFILL_17_1 gnd vdd FILL
XCLKBUF1_5 clock gnd CLKBUF1_5/Y vdd CLKBUF1
XDFFPOSX1_60 XOR2X1_3/A CLKBUF1_1/Y NOR2X1_15/Y gnd vdd DFFPOSX1
XDFFPOSX1_82 INVX1_36/A CLKBUF1_1/Y AOI21X1_19/Y gnd vdd DFFPOSX1
XDFFPOSX1_71 INVX1_8/A NOR2X1_84/A AOI21X1_15/Y gnd vdd DFFPOSX1
XDFFPOSX1_93 INVX2_2/A CLKBUF1_7/Y AOI21X1_9/Y gnd vdd DFFPOSX1
XFILL_15_2_0 gnd vdd FILL
XBUFX4_1 BUFX4_4/A gnd BUFX4_1/Y vdd BUFX4
XINVX4_1 INVX4_1/A gnd INVX4_1/Y vdd INVX4
XFILL_12_0_0 gnd vdd FILL
XFILL_4_1_0 gnd vdd FILL
XNAND3X1_4 XNOR2X1_3/A NAND3X1_4/B NAND3X1_4/C gnd NAND3X1_4/Y vdd NAND3X1
XNAND2X1_19 OAI21X1_37/Y NAND3X1_15/Y gnd NAND2X1_19/Y vdd NAND2X1
XNOR3X1_7 INVX2_8/A NOR3X1_7/B INVX2_9/A gnd NOR3X1_7/Y vdd NOR3X1
XFILL_5_1 gnd vdd FILL
XFILL_9_0_0 gnd vdd FILL
XOAI21X1_1 OR2X2_10/A OR2X2_10/B INVX2_15/A gnd NOR2X1_1/A vdd OAI21X1
XMUX2X1_5 MUX2X1_5/A MUX2X1_5/B MUX2X1_9/S gnd MUX2X1_5/Y vdd MUX2X1
XXOR2X1_4 XOR2X1_4/A INVX1_8/A gnd XOR2X1_4/Y vdd XOR2X1
XFILL_17_2 gnd vdd FILL
XCLKBUF1_6 clock gnd CLKBUF1_6/Y vdd CLKBUF1
XFILL_15_2_1 gnd vdd FILL
XDFFPOSX1_83 INVX2_5/A CLKBUF1_3/Y AOI21X1_20/Y gnd vdd DFFPOSX1
XDFFPOSX1_61 MUX2X1_5/B CLKBUF1_3/Y NOR2X1_16/Y gnd vdd DFFPOSX1
XDFFPOSX1_72 INVX2_3/A NOR2X1_75/A AOI21X1_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_50 NOR2X1_99/A CLKBUF1_8/Y NOR2X1_21/Y gnd vdd DFFPOSX1
XDFFPOSX1_94 INVX1_7/A CLKBUF1_8/Y AOI21X1_10/Y gnd vdd DFFPOSX1
XBUFX4_2 BUFX4_4/A gnd BUFX4_2/Y vdd BUFX4
XFILL_4_1_1 gnd vdd FILL
XFILL_12_0_1 gnd vdd FILL
XNAND3X1_5 NOR2X1_31/Y NOR2X1_35/Y NOR2X1_30/Y gnd NAND3X1_7/A vdd NAND3X1
XNOR3X1_8 INVX2_9/A NOR3X1_8/B NOR3X1_8/C gnd NOR3X1_8/Y vdd NOR3X1
XFILL_5_2 gnd vdd FILL
XBUFX2_50 BUFX2_50/A gnd BUFX2_50/Y vdd BUFX2
XFILL_9_0_1 gnd vdd FILL
XOAI21X1_2 OAI21X1_2/A OAI21X1_2/B INVX2_15/A gnd NOR2X1_2/A vdd OAI21X1
XXOR2X1_5 XOR2X1_5/A XOR2X1_5/B gnd XOR2X1_5/Y vdd XOR2X1
XMUX2X1_6 MUX2X1_6/A MUX2X1_6/B MUX2X1_9/S gnd MUX2X1_6/Y vdd MUX2X1
XCLKBUF1_7 clock gnd CLKBUF1_7/Y vdd CLKBUF1
XDFFPOSX1_73 INVX2_6/A NOR2X1_18/A AOI21X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_84 XOR2X1_1/B CLKBUF1_3/Y AOI21X1_21/Y gnd vdd DFFPOSX1
XDFFPOSX1_40 XOR2X1_1/A INVX8_2/A NOR2X1_27/Y gnd vdd DFFPOSX1
XDFFPOSX1_62 MUX2X1_6/B CLKBUF1_7/Y NOR2X1_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_51 XOR2X1_8/A CLKBUF1_8/Y NOR2X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_95 XOR2X1_8/B CLKBUF1_8/Y AOI21X1_11/Y gnd vdd DFFPOSX1
XBUFX4_3 BUFX4_4/A gnd BUFX4_3/Y vdd BUFX4
XNAND3X1_6 NOR2X1_31/Y NOR2X1_36/Y NOR2X1_30/Y gnd XNOR2X1_4/A vdd NAND3X1
XNOR3X1_9 XOR2X1_1/Y XOR2X1_2/Y NOR3X1_9/C gnd NOR3X1_9/Y vdd NOR3X1
XBUFX2_40 gnd gnd BUFX2_40/Y vdd BUFX2
XBUFX2_51 gnd gnd BUFX2_51/Y vdd BUFX2
XAOI21X1_30 AOI21X1_30/A NOR3X1_5/Y NOR3X1_8/Y gnd AOI21X1_31/B vdd AOI21X1
XOAI21X1_3 INVX2_1/Y INVX1_1/A INVX2_15/A gnd NOR2X1_4/B vdd OAI21X1
XMUX2X1_7 MUX2X1_7/A XOR2X1_6/A MUX2X1_9/S gnd MUX2X1_7/Y vdd MUX2X1
XFILL_10_1_0 gnd vdd FILL
XXOR2X1_6 XOR2X1_6/A INVX2_7/A gnd XOR2X1_6/Y vdd XOR2X1
XFILL_2_2_0 gnd vdd FILL
XCLKBUF1_8 clock gnd CLKBUF1_8/Y vdd CLKBUF1
XDFFPOSX1_85 INVX1_41/A CLKBUF1_2/Y AOI21X1_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_63 XOR2X1_6/A CLKBUF1_3/Y NOR2X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_74 INVX1_48/A NOR2X1_18/A AOI21X1_23/Y gnd vdd DFFPOSX1
XDFFPOSX1_41 MUX2X1_1/B NOR2X1_75/A NOR2X1_12/Y gnd vdd DFFPOSX1
XDFFPOSX1_30 AOI21X1_8/C CLKBUF1_7/Y NOR2X1_10/Y gnd vdd DFFPOSX1
XDFFPOSX1_96 INVX1_9/A CLKBUF1_7/Y NOR2X1_33/Y gnd vdd DFFPOSX1
XDFFPOSX1_52 XOR2X1_7/A CLKBUF1_8/Y NOR2X1_23/Y gnd vdd DFFPOSX1
XFILL_15_1 gnd vdd FILL
XFILL_15_0_0 gnd vdd FILL
XFILL_7_1_0 gnd vdd FILL
XBUFX4_4 BUFX4_4/A gnd BUFX4_4/Y vdd BUFX4
XNAND3X1_7 NAND3X1_7/A XNOR2X1_4/A NAND3X1_7/C gnd NAND3X1_7/Y vdd NAND3X1
XBUFX2_1 BUFX2_1/A gnd alarm_sound vdd BUFX2
XBUFX2_41 gnd gnd BUFX2_41/Y vdd BUFX2
XINVX2_1 INVX2_1/A gnd INVX2_1/Y vdd INVX2
XAOI21X1_1 AOI21X1_2/A INVX2_17/Y AOI21X1_1/C gnd AOI21X1_1/Y vdd AOI21X1
XBUFX2_52 INVX1_27/Y gnd BUFX2_52/Y vdd BUFX2
XBUFX2_30 vdd gnd ms_minute[4] vdd BUFX2
XAOI21X1_20 BUFX4_11/Y OAI21X1_29/Y OAI21X1_30/Y gnd AOI21X1_20/Y vdd AOI21X1
XOAI21X1_4 NOR2X1_4/A OAI21X1_4/B INVX2_15/A gnd OAI21X1_4/Y vdd OAI21X1
XAOI21X1_31 AOI22X1_2/Y AOI21X1_31/B NOR2X1_104/A gnd AOI21X1_31/Y vdd AOI21X1
XFILL_3_1 gnd vdd FILL
XFILL_10_1_1 gnd vdd FILL
XMUX2X1_8 MUX2X1_8/A XOR2X1_5/A MUX2X1_9/S gnd MUX2X1_8/Y vdd MUX2X1
XFILL_2_2_1 gnd vdd FILL
XXOR2X1_7 XOR2X1_7/A INVX1_9/A gnd XOR2X1_7/Y vdd XOR2X1
XCLKBUF1_9 reset gnd NOR2X1_25/A vdd CLKBUF1
XDFFPOSX1_53 NOR2X1_86/A CLKBUF1_1/Y NOR2X1_24/Y gnd vdd DFFPOSX1
XDFFPOSX1_75 INVX2_7/A NOR2X1_79/A AOI21X1_24/Y gnd vdd DFFPOSX1
XDFFPOSX1_86 INVX2_4/A CLKBUF1_2/Y NOR2X1_34/Y gnd vdd DFFPOSX1
XDFFPOSX1_42 MUX2X1_2/B NOR2X1_84/A NOR2X1_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_31 AND2X2_2/B CLKBUF1_7/Y NOR2X1_11/Y gnd vdd DFFPOSX1
XDFFPOSX1_20 AOI21X1_2/A CLKBUF1_4/Y AOI21X1_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_97 INVX1_20/A INVX2_11/A NOR2X1_52/Y gnd vdd DFFPOSX1
XDFFPOSX1_64 XOR2X1_5/A CLKBUF1_8/Y NOR2X1_19/Y gnd vdd DFFPOSX1
XFILL_15_2 gnd vdd FILL
XFILL_15_0_1 gnd vdd FILL
XFILL_7_1_1 gnd vdd FILL
XBUFX4_5 BUFX4_9/A gnd BUFX4_5/Y vdd BUFX4
XBUFX2_2 BUFX2_2/A gnd ls_hour[0] vdd BUFX2
XNAND3X1_8 INVX2_6/Y INVX1_48/A NOR2X1_37/Y gnd NOR2X1_38/B vdd NAND3X1
XINVX2_2 INVX2_2/A gnd INVX2_2/Y vdd INVX2
XAOI21X1_2 AOI21X1_2/A INVX2_17/Y AOI21X1_2/C gnd NOR2X1_1/B vdd AOI21X1
XBUFX2_31 vdd gnd ms_minute[5] vdd BUFX2
XBUFX2_20 BUFX2_20/A gnd ms_hour[2] vdd BUFX2
XBUFX2_42 vdd gnd BUFX2_42/Y vdd BUFX2
XBUFX2_53 INVX1_33/A gnd BUFX2_53/Y vdd BUFX2
XAOI21X1_21 BUFX4_12/Y NAND3X1_10/Y OAI21X1_32/Y gnd AOI21X1_21/Y vdd AOI21X1
XOAI21X1_5 OR2X2_10/Y OAI21X1_5/B INVX2_15/A gnd NOR2X1_5/A vdd OAI21X1
XAOI21X1_32 AOI22X1_4/Y AOI22X1_3/Y NOR2X1_23/A gnd AOI21X1_32/Y vdd AOI21X1
XAOI21X1_10 BUFX4_14/Y NAND3X1_3/Y OAI21X1_13/Y gnd AOI21X1_10/Y vdd AOI21X1
XFILL_3_2 gnd vdd FILL
XMUX2X1_9 MUX2X1_9/A MUX2X1_9/B MUX2X1_9/S gnd MUX2X1_9/Y vdd MUX2X1
XXOR2X1_8 XOR2X1_8/A XOR2X1_8/B gnd XOR2X1_8/Y vdd XOR2X1
XDFFPOSX1_65 INVX4_1/A NOR2X1_79/A AOI21X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_87 INVX1_8/A CLKBUF1_5/Y AOI21X1_15/Y gnd vdd DFFPOSX1
XDFFPOSX1_76 XOR2X1_5/B NOR2X1_18/A AOI21X1_25/Y gnd vdd DFFPOSX1
XDFFPOSX1_43 XOR2X1_4/A NOR2X1_75/A NOR2X1_14/Y gnd vdd DFFPOSX1
XDFFPOSX1_21 AOI21X1_2/C CLKBUF1_4/Y NOR2X1_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_10 AOI21X1_4/C NOR2X1_104/A NOR2X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_32 INVX1_59/A CLKBUF1_6/Y NOR2X1_107/Y gnd vdd DFFPOSX1
XDFFPOSX1_54 NOR2X1_87/A CLKBUF1_8/Y NOR2X1_25/Y gnd vdd DFFPOSX1
XDFFPOSX1_98 INVX1_21/A INVX2_11/A NOR2X1_53/Y gnd vdd DFFPOSX1
XNOR3X1_10 XOR2X1_3/Y XOR2X1_4/Y OAI22X1_2/Y gnd NOR3X1_10/Y vdd NOR3X1
XBUFX4_6 BUFX4_9/A gnd BUFX4_6/Y vdd BUFX4
XBUFX2_3 BUFX2_3/A gnd ls_hour[1] vdd BUFX2
XNAND3X1_9 XOR2X1_1/B INVX1_14/Y NOR2X1_41/Y gnd NAND3X1_9/Y vdd NAND3X1
XINVX2_3 INVX2_3/A gnd INVX2_3/Y vdd INVX2
XAOI21X1_3 AOI21X1_4/A INVX2_1/Y OAI21X1_4/Y gnd AOI21X1_3/Y vdd AOI21X1
XBUFX2_43 vdd gnd BUFX2_43/Y vdd BUFX2
XBUFX2_21 INVX1_51/Y gnd ms_hour[3] vdd BUFX2
XBUFX2_10 BUFX2_10/A gnd ls_minute[0] vdd BUFX2
XNOR2X1_1 NOR2X1_1/A NOR2X1_1/B gnd NOR2X1_1/Y vdd NOR2X1
XBUFX2_32 gnd gnd ms_minute[6] vdd BUFX2
XBUFX2_54 INVX1_32/A gnd BUFX2_54/Y vdd BUFX2
XAOI21X1_33 MUX2X1_35/Y NOR2X1_89/A INVX1_39/A gnd NOR2X1_88/B vdd AOI21X1
XAOI21X1_22 BUFX4_11/Y XNOR2X1_4/Y OAI21X1_33/Y gnd AOI21X1_22/Y vdd AOI21X1
XOAI21X1_6 OR2X2_1/A INVX1_4/A INVX2_15/A gnd OAI21X1_6/Y vdd OAI21X1
XFILL_5_2_0 gnd vdd FILL
XAOI21X1_11 BUFX4_14/Y NAND3X1_4/Y OAI21X1_15/Y gnd AOI21X1_11/Y vdd AOI21X1
XFILL_13_1_0 gnd vdd FILL
XDFFPOSX1_11 INVX1_2/A NOR2X1_23/A AND2X2_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_44 XOR2X1_3/A NOR2X1_77/A NOR2X1_15/Y gnd vdd DFFPOSX1
XDFFPOSX1_66 INVX1_36/A NOR2X1_84/A AOI21X1_19/Y gnd vdd DFFPOSX1
XDFFPOSX1_99 INVX2_12/A NOR2X1_75/A NOR2X1_54/Y gnd vdd DFFPOSX1
XDFFPOSX1_88 INVX2_3/A CLKBUF1_2/Y AOI21X1_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_55 XOR2X1_2/A CLKBUF1_5/Y NOR2X1_26/Y gnd vdd DFFPOSX1
XDFFPOSX1_22 OAI21X1_2/B CLKBUF1_6/Y NOR2X1_2/Y gnd vdd DFFPOSX1
XDFFPOSX1_77 INVX2_2/A NOR2X1_25/A AOI21X1_9/Y gnd vdd DFFPOSX1
XFILL_2_0_0 gnd vdd FILL
XDFFPOSX1_33 MUX2X1_9/B NOR2X1_25/A NOR2X1_20/Y gnd vdd DFFPOSX1
XNOR3X1_11 XOR2X1_5/Y XOR2X1_6/Y OAI22X1_3/Y gnd NOR3X1_11/Y vdd NOR3X1
XBUFX4_7 BUFX4_9/A gnd BUFX4_7/Y vdd BUFX4
XBUFX2_4 BUFX2_4/A gnd ls_hour[2] vdd BUFX2
XINVX2_4 INVX2_4/A gnd INVX2_4/Y vdd INVX2
XAOI21X1_4 AOI21X1_4/A INVX2_1/Y AOI21X1_4/C gnd NOR2X1_5/B vdd AOI21X1
XBUFX2_22 vdd gnd ms_hour[4] vdd BUFX2
XBUFX2_11 BUFX2_11/A gnd ls_minute[1] vdd BUFX2
XBUFX2_33 gnd gnd ms_minute[7] vdd BUFX2
XNOR2X1_2 NOR2X1_2/A INVX2_1/Y gnd NOR2X1_2/Y vdd NOR2X1
XBUFX2_44 gnd gnd BUFX2_44/Y vdd BUFX2
XBUFX2_55 OR2X2_9/B gnd BUFX2_55/Y vdd BUFX2
XAOI21X1_23 BUFX4_11/Y NAND3X1_13/Y OAI21X1_35/Y gnd AOI21X1_23/Y vdd AOI21X1
XAOI21X1_34 MUX2X1_39/Y NOR2X1_93/A INVX1_45/A gnd NOR2X1_92/B vdd AOI21X1
XOAI21X1_7 INVX1_5/Y NOR3X1_2/C INVX2_15/A gnd NOR3X1_1/A vdd OAI21X1
XAOI21X1_12 INVX1_9/A NAND3X1_4/C OAI21X1_16/Y gnd NOR2X1_33/B vdd AOI21X1
XFILL_13_1_1 gnd vdd FILL
XFILL_5_2_1 gnd vdd FILL
XFILL_1_1 gnd vdd FILL
XDFFPOSX1_67 INVX2_5/A NOR2X1_79/A AOI21X1_20/Y gnd vdd DFFPOSX1
XDFFPOSX1_89 INVX2_6/A CLKBUF1_3/Y AOI21X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_45 MUX2X1_5/B NOR2X1_18/A NOR2X1_16/Y gnd vdd DFFPOSX1
XDFFPOSX1_56 XOR2X1_1/A CLKBUF1_8/Y NOR2X1_27/Y gnd vdd DFFPOSX1
XDFFPOSX1_23 INVX1_1/A CLKBUF1_6/Y NOR2X1_4/Y gnd vdd DFFPOSX1
XFILL_2_0_1 gnd vdd FILL
XDFFPOSX1_12 INVX1_3/A NOR2X1_23/A AOI21X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_34 NOR2X1_99/A NOR2X1_23/A NOR2X1_21/Y gnd vdd DFFPOSX1
XDFFPOSX1_78 INVX1_7/A NOR2X1_25/A AOI21X1_10/Y gnd vdd DFFPOSX1
XBUFX4_8 BUFX4_9/A gnd BUFX4_8/Y vdd BUFX4
XNOR3X1_12 XOR2X1_7/Y XOR2X1_8/Y OAI22X1_4/Y gnd NOR3X1_12/Y vdd NOR3X1
XBUFX2_5 BUFX2_5/A gnd ls_hour[3] vdd BUFX2
XINVX2_5 INVX2_5/A gnd INVX2_5/Y vdd INVX2
XBUFX2_45 gnd gnd BUFX2_45/Y vdd BUFX2
XBUFX2_12 BUFX2_12/A gnd ls_minute[2] vdd BUFX2
XAOI21X1_5 OR2X2_1/B OR2X2_1/A INVX2_15/Y gnd AND2X2_1/B vdd AOI21X1
XBUFX2_34 vdd gnd BUFX2_34/Y vdd BUFX2
XBUFX2_56 BUFX2_56/A gnd BUFX2_56/Y vdd BUFX2
XBUFX2_23 vdd gnd ms_hour[5] vdd BUFX2
XAOI21X1_35 MUX2X1_43/Y NOR2X1_97/A INVX1_51/A gnd NOR2X1_96/B vdd AOI21X1
XAOI21X1_24 BUFX4_11/Y XNOR2X1_5/Y OAI21X1_36/Y gnd AOI21X1_24/Y vdd AOI21X1
XAOI21X1_13 BUFX4_13/Y XNOR2X1_2/Y OAI21X1_18/Y gnd AOI21X1_13/Y vdd AOI21X1
XNOR2X1_3 INVX1_1/Y INVX2_1/A gnd NOR2X1_4/A vdd NOR2X1
XOAI21X1_8 INVX1_6/Y OAI21X1_9/B OAI21X1_9/C gnd NOR2X1_9/B vdd OAI21X1
XFILL_1_2 gnd vdd FILL
XDFFPOSX1_57 MUX2X1_1/B CLKBUF1_2/Y NOR2X1_12/Y gnd vdd DFFPOSX1
XDFFPOSX1_68 XOR2X1_1/B NOR2X1_18/A AOI21X1_21/Y gnd vdd DFFPOSX1
XDFFPOSX1_24 OAI21X1_4/B CLKBUF1_6/Y AOI21X1_3/Y gnd vdd DFFPOSX1
XDFFPOSX1_13 NOR2X1_6/A NOR2X1_25/A NOR3X1_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_46 MUX2X1_6/B NOR2X1_25/A NOR2X1_17/Y gnd vdd DFFPOSX1
XDFFPOSX1_35 XOR2X1_8/A NOR2X1_25/A NOR2X1_22/Y gnd vdd DFFPOSX1
XDFFPOSX1_79 XOR2X1_8/B INVX8_2/A AOI21X1_11/Y gnd vdd DFFPOSX1
XFILL_11_2_0 gnd vdd FILL
XBUFX4_9 BUFX4_9/A gnd BUFX4_9/Y vdd BUFX4
XNOR3X1_13 OAI21X1_5/B INVX1_4/A OR2X2_10/Y gnd NOR2X1_6/B vdd NOR3X1
XBUFX2_6 vdd gnd ls_hour[4] vdd BUFX2
XNOR2X1_90 MUX2X1_1/B INVX1_41/A gnd OAI22X1_2/B vdd NOR2X1
XNAND2X1_1 OAI21X1_2/B OAI21X1_2/A gnd INVX2_1/A vdd NAND2X1
XFILL_16_1_0 gnd vdd FILL
XBUFX2_13 INVX1_45/Y gnd ls_minute[3] vdd BUFX2
XINVX2_6 INVX2_6/A gnd INVX2_6/Y vdd INVX2
XBUFX2_35 vdd gnd BUFX2_35/Y vdd BUFX2
XFILL_8_2_0 gnd vdd FILL
XFILL_0_1_0 gnd vdd FILL
XAOI21X1_6 INVX1_3/Y OR2X2_1/Y OAI21X1_6/Y gnd AOI21X1_6/Y vdd AOI21X1
XDFFPOSX1_1 INVX2_10/A INVX2_11/A NOR2X1_105/Y gnd vdd DFFPOSX1
XBUFX2_24 gnd gnd ms_hour[6] vdd BUFX2
XBUFX2_46 vdd gnd BUFX2_46/Y vdd BUFX2
XNOR2X1_4 NOR2X1_4/A NOR2X1_4/B gnd NOR2X1_4/Y vdd NOR2X1
XAOI21X1_36 MUX2X1_47/Y MUX2X1_48/Y INVX1_57/A gnd NOR2X1_100/B vdd AOI21X1
XAOI21X1_14 NOR2X1_30/A NOR2X1_29/Y OAI21X1_19/Y gnd NOR2X1_34/B vdd AOI21X1
XAOI21X1_25 BUFX4_12/Y NAND2X1_19/Y OAI21X1_38/Y gnd AOI21X1_25/Y vdd AOI21X1
XOAI21X1_9 NOR3X1_2/B OAI21X1_9/B OAI21X1_9/C gnd OAI21X1_9/Y vdd OAI21X1
XFILL_5_0_0 gnd vdd FILL
XDFFPOSX1_69 INVX1_41/A NOR2X1_75/A AOI21X1_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_47 XOR2X1_6/A NOR2X1_18/A NOR2X1_18/Y gnd vdd DFFPOSX1
XDFFPOSX1_58 MUX2X1_2/B CLKBUF1_1/Y NOR2X1_13/Y gnd vdd DFFPOSX1
XDFFPOSX1_14 INVX1_6/A NOR2X1_23/A NOR2X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_25 AOI21X1_4/C CLKBUF1_6/Y NOR2X1_5/Y gnd vdd DFFPOSX1
XDFFPOSX1_36 XOR2X1_7/A NOR2X1_23/A NOR2X1_23/Y gnd vdd DFFPOSX1
XFILL_11_2_1 gnd vdd FILL
XBUFX2_7 vdd gnd ls_hour[5] vdd BUFX2
XFILL_11_1 gnd vdd FILL
XNOR2X1_91 MUX2X1_2/B INVX2_4/A gnd OAI22X1_2/D vdd NOR2X1
XNOR2X1_80 INVX8_2/A NOR2X1_80/B gnd NOR2X1_80/Y vdd NOR2X1
XINVX2_7 INVX2_7/A gnd INVX2_7/Y vdd INVX2
XINVX1_50 XOR2X1_5/B gnd INVX1_50/Y vdd INVX1
XFILL_8_2_1 gnd vdd FILL
XFILL_0_1_1 gnd vdd FILL
XAOI21X1_7 INVX1_5/A NOR2X1_6/B INVX2_15/Y gnd OAI21X1_9/C vdd AOI21X1
XNAND2X1_2 NOR2X1_6/A NOR2X1_6/B gnd OAI21X1_9/B vdd NAND2X1
XBUFX2_14 vdd gnd ls_minute[4] vdd BUFX2
XFILL_16_1_1 gnd vdd FILL
XNOR2X1_5 NOR2X1_5/A NOR2X1_5/B gnd NOR2X1_5/Y vdd NOR2X1
XDFFPOSX1_2 INVX2_10/A CLKBUF1_4/Y NOR2X1_105/Y gnd vdd DFFPOSX1
XBUFX2_47 vdd gnd BUFX2_47/Y vdd BUFX2
XBUFX2_36 gnd gnd BUFX2_36/Y vdd BUFX2
XBUFX2_25 gnd gnd ms_hour[7] vdd BUFX2
XAOI21X1_15 BUFX4_10/Y NAND2X1_12/Y OAI21X1_22/Y gnd AOI21X1_15/Y vdd AOI21X1
XAOI21X1_26 OAI21X1_42/Y NAND2X1_26/Y NOR2X1_53/B gnd AOI21X1_26/Y vdd AOI21X1
XFILL_5_0_1 gnd vdd FILL
XDFFPOSX1_37 NOR2X1_86/A NOR2X1_77/A NOR2X1_24/Y gnd vdd DFFPOSX1
XDFFPOSX1_59 XOR2X1_4/A CLKBUF1_5/Y NOR2X1_14/Y gnd vdd DFFPOSX1
XDFFPOSX1_26 INVX1_2/A CLKBUF1_7/Y AND2X2_1/Y gnd vdd DFFPOSX1
XDFFPOSX1_15 AOI21X1_8/C NOR2X1_25/A NOR2X1_10/Y gnd vdd DFFPOSX1
XDFFPOSX1_48 XOR2X1_5/A NOR2X1_18/A NOR2X1_19/Y gnd vdd DFFPOSX1
XBUFX2_8 gnd gnd ls_hour[6] vdd BUFX2
XNOR2X1_70 NOR2X1_79/A NOR2X1_70/B gnd NOR2X1_70/Y vdd NOR2X1
XNOR2X1_92 NOR2X1_92/A NOR2X1_92/B gnd BUFX2_10/A vdd NOR2X1
XNOR2X1_81 INVX8_2/A NOR2X1_81/B gnd NOR2X1_81/Y vdd NOR2X1
XNAND2X1_3 INVX1_41/A XNOR2X1_2/B gnd INVX1_11/A vdd NAND2X1
XAOI21X1_8 INVX1_6/A NOR3X1_1/B AOI21X1_8/C gnd NOR2X1_10/A vdd AOI21X1
XINVX2_8 INVX2_8/A gnd INVX2_8/Y vdd INVX2
XBUFX2_15 vdd gnd ls_minute[5] vdd BUFX2
XBUFX2_26 BUFX2_26/A gnd ms_minute[0] vdd BUFX2
XINVX1_51 INVX1_51/A gnd INVX1_51/Y vdd INVX1
XINVX1_40 BUFX4_1/Y gnd INVX1_40/Y vdd INVX1
XBUFX2_37 gnd gnd BUFX2_37/Y vdd BUFX2
XNOR2X1_6 NOR2X1_6/A NOR2X1_6/B gnd NOR3X1_1/C vdd NOR2X1
XDFFPOSX1_3 OAI21X1_67/A INVX2_11/A NOR2X1_108/Y gnd vdd DFFPOSX1
XBUFX2_48 gnd gnd BUFX2_48/Y vdd BUFX2
XAOI21X1_16 INVX2_3/Y OR2X2_3/Y NOR2X1_30/Y gnd OAI21X1_23/C vdd AOI21X1
XAOI21X1_27 OAI21X1_45/Y NAND2X1_29/Y NOR2X1_60/B gnd AOI21X1_27/Y vdd AOI21X1
XDFFPOSX1_16 AND2X2_2/B NOR2X1_23/A NOR2X1_11/Y gnd vdd DFFPOSX1
XDFFPOSX1_27 INVX1_3/A CLKBUF1_6/Y AOI21X1_6/Y gnd vdd DFFPOSX1
XDFFPOSX1_49 MUX2X1_9/B CLKBUF1_7/Y NOR2X1_20/Y gnd vdd DFFPOSX1
XDFFPOSX1_38 NOR2X1_87/A NOR2X1_18/A NOR2X1_25/Y gnd vdd DFFPOSX1
XFILL_14_2_0 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XNOR2X1_71 NOR2X1_79/A NOR2X1_71/B gnd NOR2X1_71/Y vdd NOR2X1
XNOR2X1_93 NOR2X1_93/A INVX1_45/Y gnd BUFX2_12/A vdd NOR2X1
XFILL_11_0_0 gnd vdd FILL
XNOR2X1_82 NOR2X1_84/A NOR2X1_82/B gnd NOR2X1_82/Y vdd NOR2X1
XNOR2X1_60 NOR2X1_60/A NOR2X1_60/B gnd NOR2X1_60/Y vdd NOR2X1
XBUFX2_9 gnd gnd ls_hour[7] vdd BUFX2
XNAND2X1_4 NOR2X1_28/Y NOR2X1_29/Y gnd OR2X2_2/A vdd NAND2X1
XAOI21X1_9 BUFX4_12/Y XNOR2X1_1/Y AOI21X1_9/C gnd AOI21X1_9/Y vdd AOI21X1
XINVX2_9 INVX2_9/A gnd OR2X2_9/A vdd INVX2
XBUFX2_16 gnd gnd ls_minute[6] vdd BUFX2
XBUFX2_27 BUFX2_27/A gnd ms_minute[1] vdd BUFX2
XINVX1_52 BUFX4_4/Y gnd INVX1_52/Y vdd INVX1
XINVX1_41 INVX1_41/A gnd INVX1_41/Y vdd INVX1
XBUFX2_49 gnd gnd BUFX2_49/Y vdd BUFX2
XNOR2X1_7 NOR3X1_2/A NOR3X1_2/C gnd NOR3X1_1/B vdd NOR2X1
XINVX1_30 INVX1_30/A gnd INVX1_30/Y vdd INVX1
XDFFPOSX1_4 OAI21X1_67/B INVX2_11/A NOR2X1_109/Y gnd vdd DFFPOSX1
XBUFX2_38 vdd gnd BUFX2_38/Y vdd BUFX2
XAOI21X1_17 BUFX4_13/Y OAI21X1_23/Y OAI21X1_24/Y gnd AOI21X1_17/Y vdd AOI21X1
XAOI21X1_28 AOI21X1_28/A NOR3X1_6/Y NOR3X1_8/Y gnd AOI21X1_29/B vdd AOI21X1
XFILL_8_0_0 gnd vdd FILL
XDFFPOSX1_39 XOR2X1_2/A NOR2X1_84/A NOR2X1_26/Y gnd vdd DFFPOSX1
XDFFPOSX1_17 INVX1_59/A NOR2X1_104/A NOR2X1_107/Y gnd vdd DFFPOSX1
XDFFPOSX1_28 NOR2X1_6/A CLKBUF1_7/Y NOR3X1_1/Y gnd vdd DFFPOSX1
XFILL_14_2_1 gnd vdd FILL
XFILL_3_1_1 gnd vdd FILL
XNOR2X1_72 NOR2X1_79/A NOR2X1_72/B gnd NOR2X1_72/Y vdd NOR2X1
XFILL_11_0_1 gnd vdd FILL
XNOR2X1_94 MUX2X1_5/B INVX2_6/A gnd OAI22X1_3/B vdd NOR2X1
XNOR2X1_83 INVX8_2/A NOR2X1_83/B gnd NOR2X1_83/Y vdd NOR2X1
XNOR2X1_50 INVX2_10/A INVX1_20/Y gnd NOR2X1_50/Y vdd NOR2X1
XNOR2X1_61 NOR2X1_61/A XNOR2X1_7/Y gnd NOR2X1_61/Y vdd NOR2X1
XNAND2X1_5 INVX2_2/A INVX1_7/A gnd OR2X2_2/B vdd NAND2X1
XBUFX2_28 BUFX2_28/A gnd ms_minute[2] vdd BUFX2
XINVX1_42 INVX2_4/A gnd INVX1_42/Y vdd INVX1
XINVX1_20 INVX1_20/A gnd INVX1_20/Y vdd INVX1
XBUFX2_17 gnd gnd ls_minute[7] vdd BUFX2
XINVX1_31 time_button gnd INVX1_31/Y vdd INVX1
XDFFPOSX1_5 AOI21X1_2/A INVX2_11/A AOI21X1_1/Y gnd vdd DFFPOSX1
XBUFX2_39 vdd gnd BUFX2_39/Y vdd BUFX2
XINVX1_53 INVX2_2/A gnd INVX1_53/Y vdd INVX1
XAOI21X1_18 BUFX4_10/Y XNOR2X1_3/Y OAI21X1_25/Y gnd AOI21X1_18/Y vdd AOI21X1
XNOR2X1_8 INVX1_6/A NOR3X1_1/B gnd NOR2X1_9/A vdd NOR2X1
XAOI21X1_29 AOI22X1_1/Y AOI21X1_29/B NOR2X1_104/A gnd AOI21X1_29/Y vdd AOI21X1
XFILL_8_0_1 gnd vdd FILL
XDFFPOSX1_29 INVX1_6/A CLKBUF1_7/Y NOR2X1_9/Y gnd vdd DFFPOSX1
XDFFPOSX1_18 OAI21X1_67/A CLKBUF1_4/Y NOR2X1_108/Y gnd vdd DFFPOSX1
XNOR2X1_73 NOR2X1_77/A NOR2X1_73/B gnd NOR2X1_73/Y vdd NOR2X1
XNAND2X1_6 INVX2_3/A OR2X2_3/B gnd NOR2X1_30/A vdd NAND2X1
XNOR2X1_95 MUX2X1_6/B INVX1_48/A gnd OAI22X1_3/D vdd NOR2X1
XNOR2X1_84 NOR2X1_84/A NOR2X1_84/B gnd NOR2X1_84/Y vdd NOR2X1
XNOR2X1_62 INVX2_13/Y XNOR2X1_7/A gnd NOR2X1_62/Y vdd NOR2X1
XNOR2X1_51 INVX1_20/A INVX2_10/Y gnd NOR2X1_51/Y vdd NOR2X1
XNOR2X1_40 INVX1_9/A INVX1_10/Y gnd NOR2X1_40/Y vdd NOR2X1
XBUFX2_29 INVX1_57/Y gnd ms_minute[3] vdd BUFX2
XBUFX2_18 BUFX2_18/A gnd ms_hour[0] vdd BUFX2
XINVX1_43 INVX1_8/A gnd INVX1_43/Y vdd INVX1
XINVX1_21 INVX1_21/A gnd INVX1_21/Y vdd INVX1
XDFFPOSX1_6 AOI21X1_2/C INVX2_11/A NOR2X1_1/Y gnd vdd DFFPOSX1
XINVX1_32 INVX1_32/A gnd INVX1_32/Y vdd INVX1
XINVX1_54 INVX1_7/A gnd INVX1_54/Y vdd INVX1
XINVX1_10 XOR2X1_8/B gnd INVX1_10/Y vdd INVX1
XNOR2X1_9 NOR2X1_9/A NOR2X1_9/B gnd NOR2X1_9/Y vdd NOR2X1
XAOI21X1_19 BUFX4_10/Y NAND3X1_7/Y OAI21X1_27/Y gnd AOI21X1_19/Y vdd AOI21X1
XOAI21X1_60 INVX1_51/A NOR2X1_97/A MUX2X1_43/Y gnd BUFX2_19/A vdd OAI21X1
XFILL_8_1 gnd vdd FILL
XFILL_1_2_0 gnd vdd FILL
XDFFPOSX1_19 OAI21X1_67/B CLKBUF1_4/Y NOR2X1_109/Y gnd vdd DFFPOSX1
XFILL_14_0_0 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XNOR2X1_74 NOR2X1_75/A NOR2X1_74/B gnd NOR2X1_74/Y vdd NOR2X1
XNOR2X1_96 NOR2X1_96/A NOR2X1_96/B gnd BUFX2_18/A vdd NOR2X1
XNOR2X1_30 NOR2X1_30/A NOR2X1_30/B gnd NOR2X1_30/Y vdd NOR2X1
XNOR2X1_41 NOR3X1_4/B OR2X2_2/A gnd NOR2X1_41/Y vdd NOR2X1
XNOR2X1_85 NOR2X1_85/A NOR2X1_85/B gnd BUFX2_1/A vdd NOR2X1
XNAND2X1_7 INVX2_2/A INVX1_7/Y gnd NOR2X1_31/A vdd NAND2X1
XNOR2X1_63 INVX1_28/Y INVX1_27/A gnd NOR2X1_63/Y vdd NOR2X1
XNOR2X1_52 NOR2X1_54/B NOR2X1_52/B gnd NOR2X1_52/Y vdd NOR2X1
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XINVX1_44 INVX2_3/A gnd INVX1_44/Y vdd INVX1
XINVX1_22 INVX1_22/A gnd INVX1_22/Y vdd INVX1
XINVX1_33 INVX1_33/A gnd NOR3X1_8/B vdd INVX1
XINVX1_55 XOR2X1_8/B gnd INVX1_55/Y vdd INVX1
XBUFX2_19 BUFX2_19/A gnd ms_hour[1] vdd BUFX2
XDFFPOSX1_7 OAI21X1_2/B NOR2X1_104/A NOR2X1_2/Y gnd vdd DFFPOSX1
XOAI21X1_50 INVX1_39/A NOR2X1_89/A MUX2X1_35/Y gnd BUFX2_3/A vdd OAI21X1
XFILL_8_2 gnd vdd FILL
XOAI21X1_61 INVX1_53/Y BUFX4_7/Y OAI21X1_61/C gnd OAI21X1_61/Y vdd OAI21X1
XFILL_1_2_1 gnd vdd FILL
XAND2X2_20 INVX1_1/A OAI21X1_4/B gnd AOI21X1_4/A vdd AND2X2
XFILL_14_0_1 gnd vdd FILL
XFILL_6_1_1 gnd vdd FILL
XNOR2X1_97 NOR2X1_97/A INVX1_51/Y gnd BUFX2_20/A vdd NOR2X1
XNOR2X1_75 NOR2X1_75/A NOR2X1_75/B gnd NOR2X1_75/Y vdd NOR2X1
XNOR2X1_42 INVX1_36/A INVX4_1/Y gnd NOR2X1_42/Y vdd NOR2X1
XNOR2X1_86 NOR2X1_86/A INVX4_1/A gnd OAI22X1_1/B vdd NOR2X1
XNOR2X1_31 NOR2X1_31/A NOR2X1_31/B gnd NOR2X1_31/Y vdd NOR2X1
XNOR2X1_53 NOR2X1_53/A NOR2X1_53/B gnd NOR2X1_53/Y vdd NOR2X1
XNOR2X1_64 INVX1_29/Y INVX1_27/A gnd NOR2X1_64/Y vdd NOR2X1
XNAND3X1_20 INVX2_10/A INVX1_23/A INVX1_24/A gnd XNOR2X1_7/A vdd NAND3X1
XNOR2X1_20 NOR2X1_25/A MUX2X1_9/Y gnd NOR2X1_20/Y vdd NOR2X1
XNAND2X1_8 XOR2X1_8/B INVX1_9/Y gnd NOR2X1_31/B vdd NAND2X1
XINVX1_12 INVX1_36/A gnd INVX1_12/Y vdd INVX1
XDFFPOSX1_8 INVX1_1/A NOR2X1_104/A NOR2X1_4/Y gnd vdd DFFPOSX1
XINVX1_23 INVX1_23/A gnd INVX1_23/Y vdd INVX1
XINVX1_34 INVX1_34/A gnd INVX1_34/Y vdd INVX1
XINVX1_56 INVX1_9/A gnd INVX1_56/Y vdd INVX1
XINVX1_45 INVX1_45/A gnd INVX1_45/Y vdd INVX1
XOAI21X1_51 INVX1_41/Y BUFX4_5/Y OAI21X1_51/C gnd OAI21X1_51/Y vdd OAI21X1
XOAI21X1_62 INVX1_54/Y BUFX4_7/Y OAI21X1_62/C gnd OAI21X1_62/Y vdd OAI21X1
XOAI21X1_40 NOR2X1_50/Y NOR2X1_51/Y OAI21X1_40/C gnd NOR2X1_52/B vdd OAI21X1
XAND2X2_10 NOR3X1_6/Y INVX1_26/A gnd AND2X2_10/Y vdd AND2X2
XNOR2X1_76 NOR2X1_77/A NOR2X1_76/B gnd NOR2X1_76/Y vdd NOR2X1
XNOR2X1_43 INVX2_5/A INVX1_13/Y gnd NOR2X1_43/Y vdd NOR2X1
XNAND3X1_10 XNOR2X1_4/A OAI21X1_31/Y NAND3X1_9/Y gnd NAND3X1_10/Y vdd NAND3X1
XNOR2X1_87 NOR2X1_87/A INVX1_36/A gnd OAI22X1_1/D vdd NOR2X1
XNOR2X1_54 XNOR2X1_6/Y NOR2X1_54/B gnd NOR2X1_54/Y vdd NOR2X1
XNOR2X1_10 NOR2X1_10/A OAI21X1_9/Y gnd NOR2X1_10/Y vdd NOR2X1
XNOR2X1_98 MUX2X1_9/B INVX2_2/A gnd OAI22X1_4/B vdd NOR2X1
XNOR2X1_65 INVX1_30/Y INVX1_27/A gnd NOR2X1_65/Y vdd NOR2X1
XNOR2X1_21 NOR2X1_23/A NOR2X1_21/B gnd NOR2X1_21/Y vdd NOR2X1
XNAND3X1_21 INVX2_11/Y NOR3X1_5/Y OAI21X1_43/C gnd NOR2X1_60/B vdd NAND3X1
XNOR2X1_32 OR2X2_2/B OR2X2_2/A gnd NOR2X1_32/Y vdd NOR2X1
XNOR2X1_100 MUX2X1_45/Y NOR2X1_100/B gnd BUFX2_26/A vdd NOR2X1
XNAND2X1_9 NOR2X1_31/Y NOR2X1_30/Y gnd XNOR2X1_3/A vdd NAND2X1
XINVX1_57 INVX1_57/A gnd INVX1_57/Y vdd INVX1
XINVX1_46 BUFX4_2/Y gnd INVX1_46/Y vdd INVX1
XINVX1_35 INVX4_1/A gnd INVX1_35/Y vdd INVX1
XINVX1_13 XOR2X1_1/B gnd INVX1_13/Y vdd INVX1
XDFFPOSX1_9 OAI21X1_4/B INVX2_11/A AOI21X1_3/Y gnd vdd DFFPOSX1
XINVX1_24 INVX1_24/A gnd INVX1_24/Y vdd INVX1
XFILL_12_1_0 gnd vdd FILL
XFILL_4_2_0 gnd vdd FILL
XOAI21X1_30 BUFX4_10/Y MUX2X1_36/A INVX8_2/Y gnd OAI21X1_30/Y vdd OAI21X1
XOAI21X1_52 INVX1_42/Y BUFX4_5/Y OAI21X1_52/C gnd OAI21X1_52/Y vdd OAI21X1
XOAI21X1_41 INVX2_10/Y INVX1_20/Y INVX1_21/Y gnd OAI21X1_41/Y vdd OAI21X1
XOAI21X1_63 INVX1_55/Y BUFX4_7/Y OAI21X1_63/C gnd OAI21X1_63/Y vdd OAI21X1
XAND2X2_11 NOR2X1_86/A INVX4_1/A gnd OAI22X1_1/A vdd AND2X2
XFILL_6_1 gnd vdd FILL
XFILL_1_0_0 gnd vdd FILL
XFILL_9_1_0 gnd vdd FILL
XNOR2X1_88 NOR2X1_88/A NOR2X1_88/B gnd BUFX2_2/A vdd NOR2X1
XNOR2X1_44 key[0] key[2] gnd NOR2X1_44/Y vdd NOR2X1
XNOR2X1_77 NOR2X1_77/A NOR2X1_77/B gnd NOR2X1_77/Y vdd NOR2X1
XNAND3X1_11 NOR2X1_30/Y NOR2X1_31/Y NOR3X1_3/Y gnd XNOR2X1_5/A vdd NAND3X1
XNOR2X1_55 INVX2_12/Y XNOR2X1_6/A gnd NOR2X1_55/Y vdd NOR2X1
XNOR2X1_11 AND2X2_2/Y NOR2X1_11/B gnd NOR2X1_11/Y vdd NOR2X1
XNAND3X1_22 INVX1_31/Y INVX2_14/Y NOR3X1_5/Y gnd INVX1_34/A vdd NAND3X1
XNOR2X1_99 NOR2X1_99/A INVX1_7/A gnd OAI22X1_4/D vdd NOR2X1
XNOR2X1_66 alarm_button INVX1_32/Y gnd NOR2X1_66/Y vdd NOR2X1
XNOR2X1_22 NOR2X1_25/A NOR2X1_22/B gnd NOR2X1_22/Y vdd NOR2X1
XNOR2X1_33 NOR2X1_33/A NOR2X1_33/B gnd NOR2X1_33/Y vdd NOR2X1
XNOR2X1_101 MUX2X1_48/Y INVX1_57/Y gnd BUFX2_28/A vdd NOR2X1
XMUX2X1_40 MUX2X1_3/A MUX2X1_40/B BUFX4_4/Y gnd NOR2X1_93/A vdd MUX2X1
XINVX1_58 BUFX4_1/Y gnd INVX1_58/Y vdd INVX1
XINVX1_14 INVX1_14/A gnd INVX1_14/Y vdd INVX1
XINVX1_36 INVX1_36/A gnd INVX1_36/Y vdd INVX1
XINVX1_47 INVX2_6/A gnd INVX1_47/Y vdd INVX1
XINVX1_25 INVX1_25/A gnd INVX1_25/Y vdd INVX1
XFILL_12_1_1 gnd vdd FILL
XFILL_4_2_1 gnd vdd FILL
XOAI21X1_20 BUFX4_13/Y MUX2X1_2/A INVX8_2/Y gnd NOR2X1_34/A vdd OAI21X1
XOAI21X1_31 XNOR2X1_3/A INVX1_14/A INVX1_13/Y gnd OAI21X1_31/Y vdd OAI21X1
XOAI21X1_53 INVX1_43/Y BUFX4_5/Y OAI21X1_53/C gnd OAI21X1_53/Y vdd OAI21X1
XOAI21X1_42 XNOR2X1_6/A INVX2_12/Y INVX1_22/A gnd OAI21X1_42/Y vdd OAI21X1
XOAI21X1_64 INVX1_56/Y BUFX4_7/Y OAI21X1_64/C gnd OAI21X1_64/Y vdd OAI21X1
XAND2X2_12 NOR2X1_87/A INVX1_36/A gnd OAI22X1_1/C vdd AND2X2
XFILL_1_0_1 gnd vdd FILL
XCLKBUF1_10 reset gnd INVX8_2/A vdd CLKBUF1
XFILL_9_1_1 gnd vdd FILL
XNAND3X1_12 NOR2X1_35/Y NOR2X1_38/Y NOR2X1_41/Y gnd NAND3X1_13/B vdd NAND3X1
XNOR2X1_12 NOR2X1_75/A MUX2X1_1/Y gnd NOR2X1_12/Y vdd NOR2X1
XNOR2X1_89 NOR2X1_89/A BUFX2_5/A gnd BUFX2_4/A vdd NOR2X1
XMUX2X1_41 MUX2X1_5/A MUX2X1_41/B BUFX4_2/Y gnd NOR2X1_96/A vdd MUX2X1
XNOR2X1_34 NOR2X1_34/A NOR2X1_34/B gnd NOR2X1_34/Y vdd NOR2X1
XMUX2X1_30 MUX2X1_2/A MUX2X1_47/A AND2X2_4/Y gnd NOR2X1_82/B vdd MUX2X1
XNOR2X1_78 NOR2X1_84/A NOR2X1_78/B gnd NOR2X1_78/Y vdd NOR2X1
XNOR2X1_102 NOR2X1_102/A NOR2X1_102/B gnd NAND3X1_1/B vdd NOR2X1
XNOR2X1_67 alarm_button INVX1_19/Y gnd NOR2X1_67/Y vdd NOR2X1
XNOR2X1_45 INVX2_9/A NOR3X1_8/C gnd BUFX4_9/A vdd NOR2X1
XNOR2X1_23 NOR2X1_23/A NOR2X1_23/B gnd NOR2X1_23/Y vdd NOR2X1
XNOR2X1_56 INVX1_24/A INVX2_13/A gnd NOR2X1_56/Y vdd NOR2X1
XINVX1_26 INVX1_26/A gnd OR2X2_7/A vdd INVX1
XINVX1_15 INVX1_48/A gnd INVX1_15/Y vdd INVX1
XINVX1_48 INVX1_48/A gnd INVX1_48/Y vdd INVX1
XINVX1_37 INVX2_5/A gnd INVX1_37/Y vdd INVX1
XINVX1_59 INVX1_59/A gnd INVX1_59/Y vdd INVX1
XOAI21X1_65 INVX1_57/A MUX2X1_48/Y MUX2X1_47/Y gnd BUFX2_27/A vdd OAI21X1
XOAI21X1_21 INVX1_11/A INVX2_4/Y OR2X2_3/B gnd OAI21X1_21/Y vdd OAI21X1
XOAI21X1_32 BUFX4_12/Y MUX2X1_34/A INVX8_2/Y gnd OAI21X1_32/Y vdd OAI21X1
XOAI21X1_54 INVX1_44/Y BUFX4_6/Y OAI21X1_54/C gnd OAI21X1_54/Y vdd OAI21X1
XOAI21X1_10 AND2X2_2/B NOR3X1_2/Y OAI21X1_9/C gnd NOR2X1_11/B vdd OAI21X1
XOAI21X1_43 NOR2X1_57/Y NOR2X1_58/Y OAI21X1_43/C gnd NOR2X1_59/B vdd OAI21X1
XAND2X2_13 MUX2X1_1/B INVX1_41/A gnd OAI22X1_2/A vdd AND2X2
XCLKBUF1_11 reset gnd NOR2X1_84/A vdd CLKBUF1
XFILL_10_2_0 gnd vdd FILL
XNOR2X1_24 NOR2X1_79/A NOR2X1_24/B gnd NOR2X1_24/Y vdd NOR2X1
XNOR2X1_79 NOR2X1_79/A NOR2X1_79/B gnd NOR2X1_79/Y vdd NOR2X1
XNAND3X1_13 XNOR2X1_5/A NAND3X1_13/B OAI21X1_34/Y gnd NAND3X1_13/Y vdd NAND3X1
XNOR2X1_35 INVX4_1/Y INVX1_12/Y gnd NOR2X1_35/Y vdd NOR2X1
XNOR2X1_13 NOR2X1_84/A MUX2X1_2/Y gnd NOR2X1_13/Y vdd NOR2X1
XNOR2X1_57 INVX1_23/A INVX2_10/Y gnd NOR2X1_57/Y vdd NOR2X1
XNOR2X1_68 INVX1_27/A INVX1_34/A gnd NOR2X1_68/Y vdd NOR2X1
XNOR2X1_46 NOR3X1_7/B INVX2_8/Y gnd AND2X2_4/A vdd NOR2X1
XFILL_16_1 gnd vdd FILL
XMUX2X1_42 MUX2X1_8/A MUX2X1_42/B BUFX4_2/Y gnd INVX1_51/A vdd MUX2X1
XMUX2X1_20 MUX2X1_34/A MUX2X1_8/A AND2X2_4/Y gnd NOR2X1_72/B vdd MUX2X1
XINVX1_16 XOR2X1_5/B gnd INVX1_16/Y vdd INVX1
XINVX1_49 INVX2_7/A gnd INVX1_49/Y vdd INVX1
XINVX1_38 XOR2X1_1/B gnd INVX1_38/Y vdd INVX1
XMUX2X1_31 MUX2X1_3/A MUX2X1_48/A AND2X2_4/Y gnd NOR2X1_83/B vdd MUX2X1
XNOR2X1_103 OR2X2_10/A OR2X2_10/B gnd OAI21X1_2/A vdd NOR2X1
XINVX1_27 INVX1_27/A gnd INVX1_27/Y vdd INVX1
XFILL_7_2_0 gnd vdd FILL
XFILL_15_1_0 gnd vdd FILL
XOAI21X1_33 BUFX4_11/Y MUX2X1_5/A INVX8_2/Y gnd OAI21X1_33/Y vdd OAI21X1
XOAI21X1_22 BUFX4_10/Y MUX2X1_3/A INVX8_2/Y gnd OAI21X1_22/Y vdd OAI21X1
XOAI21X1_55 INVX1_45/A NOR2X1_93/A MUX2X1_39/Y gnd BUFX2_11/A vdd OAI21X1
XOAI21X1_11 BUFX4_12/Y MUX2X1_9/A INVX8_2/Y gnd AOI21X1_9/C vdd OAI21X1
XOAI21X1_66 INVX1_59/Y fastwatch OAI21X1_66/C gnd XNOR2X1_2/B vdd OAI21X1
XOAI21X1_44 INVX2_10/Y INVX1_23/Y INVX1_24/Y gnd OAI21X1_44/Y vdd OAI21X1
XAND2X2_14 MUX2X1_2/B INVX2_4/A gnd OAI22X1_2/C vdd AND2X2
XDFFPOSX1_150 MUX2X1_46/A CLKBUF1_5/Y NOR2X1_84/Y gnd vdd DFFPOSX1
XFILL_4_0_0 gnd vdd FILL
XCLKBUF1_12 reset gnd NOR2X1_104/A vdd CLKBUF1
XFILL_4_1 gnd vdd FILL
XFILL_10_2_1 gnd vdd FILL
XNOR2X1_69 NOR2X1_77/A NOR2X1_69/B gnd NOR2X1_69/Y vdd NOR2X1
XNOR2X1_36 NOR3X1_3/A NOR3X1_3/C gnd NOR2X1_36/Y vdd NOR2X1
XNAND3X1_14 INVX1_17/Y NOR2X1_42/Y NOR2X1_43/Y gnd NOR3X1_4/C vdd NAND3X1
XNOR2X1_14 INVX8_2/A MUX2X1_3/Y gnd NOR2X1_14/Y vdd NOR2X1
XNOR2X1_47 OR2X2_9/A NOR2X1_47/B gnd MUX2X1_9/S vdd NOR2X1
XNOR2X1_58 INVX2_10/A INVX1_23/Y gnd NOR2X1_58/Y vdd NOR2X1
XNOR2X1_25 NOR2X1_25/A NOR2X1_25/B gnd NOR2X1_25/Y vdd NOR2X1
XMUX2X1_21 key[0] MUX2X1_1/A AND2X2_4/Y gnd NOR2X1_73/B vdd MUX2X1
XMUX2X1_43 MUX2X1_6/A MUX2X1_43/B BUFX4_2/Y gnd MUX2X1_43/Y vdd MUX2X1
XMUX2X1_32 MUX2X1_4/A MUX2X1_46/A AND2X2_4/Y gnd NOR2X1_84/B vdd MUX2X1
XNOR2X1_104 NOR2X1_104/A INVX8_1/A gnd INVX2_15/A vdd NOR2X1
XMUX2X1_10 MUX2X1_47/A NOR2X1_99/A MUX2X1_9/S gnd NOR2X1_21/B vdd MUX2X1
XINVX1_39 INVX1_39/A gnd BUFX2_5/A vdd INVX1
XINVX1_17 NOR3X1_3/B gnd INVX1_17/Y vdd INVX1
XINVX1_28 INVX1_28/A gnd INVX1_28/Y vdd INVX1
XFILL_7_2_1 gnd vdd FILL
XFILL_15_1_1 gnd vdd FILL
XOAI21X1_23 INVX2_3/Y OR2X2_3/Y OAI21X1_23/C gnd OAI21X1_23/Y vdd OAI21X1
XOAI21X1_34 XNOR2X1_4/A INVX2_6/Y INVX1_15/Y gnd OAI21X1_34/Y vdd OAI21X1
XOAI21X1_12 OR2X2_2/A INVX2_2/Y INVX1_7/Y gnd NAND3X1_3/A vdd OAI21X1
XOAI21X1_45 XNOR2X1_7/A INVX2_13/Y INVX1_25/A gnd OAI21X1_45/Y vdd OAI21X1
XOAI21X1_56 INVX1_47/Y BUFX4_9/Y OAI21X1_56/C gnd OAI21X1_56/Y vdd OAI21X1
XOAI21X1_67 OAI21X1_67/A OAI21X1_67/B INVX2_15/A gnd OAI21X1_67/Y vdd OAI21X1
XDFFPOSX1_140 MUX2X1_2/A CLKBUF1_2/Y NOR2X1_74/Y gnd vdd DFFPOSX1
XAND2X2_15 MUX2X1_5/B INVX2_6/A gnd OAI22X1_3/A vdd AND2X2
XFILL_4_0_1 gnd vdd FILL
XCLKBUF1_13 reset gnd NOR2X1_23/A vdd CLKBUF1
XFILL_4_2 gnd vdd FILL
XNOR2X1_15 NOR2X1_77/A MUX2X1_4/Y gnd NOR2X1_15/Y vdd NOR2X1
XNOR2X1_37 XOR2X1_5/B INVX2_7/A gnd NOR2X1_37/Y vdd NOR2X1
XNAND3X1_15 XOR2X1_5/B INVX2_7/A NOR3X1_4/Y gnd NAND3X1_15/Y vdd NAND3X1
XNOR2X1_26 NOR2X1_84/A NOR2X1_26/B gnd NOR2X1_26/Y vdd NOR2X1
XNOR2X1_48 OR2X2_9/A NOR2X1_48/B gnd INVX8_1/A vdd NOR2X1
XNOR2X1_59 NOR2X1_61/A NOR2X1_59/B gnd NOR2X1_59/Y vdd NOR2X1
XMUX2X1_22 key[1] MUX2X1_2/A AND2X2_4/Y gnd NOR2X1_74/B vdd MUX2X1
XMUX2X1_44 MUX2X1_7/A MUX2X1_44/B BUFX4_2/Y gnd NOR2X1_97/A vdd MUX2X1
XMUX2X1_33 MUX2X1_33/A MUX2X1_33/B BUFX4_3/Y gnd NOR2X1_88/A vdd MUX2X1
XNOR2X1_105 INVX2_15/Y OR2X2_1/A gnd NOR2X1_105/Y vdd NOR2X1
XMUX2X1_11 MUX2X1_48/A XOR2X1_8/A MUX2X1_9/S gnd NOR2X1_22/B vdd MUX2X1
XINVX1_29 INVX1_29/A gnd INVX1_29/Y vdd INVX1
XINVX1_18 NOR3X1_7/B gnd NOR3X1_5/C vdd INVX1
XOAI21X1_24 BUFX4_13/Y MUX2X1_4/A INVX8_2/Y gnd OAI21X1_24/Y vdd OAI21X1
XOAI21X1_35 BUFX4_11/Y MUX2X1_6/A INVX8_2/Y gnd OAI21X1_35/Y vdd OAI21X1
XOAI21X1_46 INVX1_35/Y BUFX4_5/Y OAI21X1_46/C gnd OAI21X1_46/Y vdd OAI21X1
XOAI21X1_57 INVX1_48/Y BUFX4_9/Y OAI21X1_57/C gnd OAI21X1_57/Y vdd OAI21X1
XOAI21X1_68 INVX2_17/Y AOI21X1_2/A INVX2_15/A gnd AOI21X1_1/C vdd OAI21X1
XOAI21X1_13 BUFX4_14/Y MUX2X1_47/A INVX8_2/Y gnd OAI21X1_13/Y vdd OAI21X1
XDFFPOSX1_141 MUX2X1_3/A CLKBUF1_2/Y NOR2X1_75/Y gnd vdd DFFPOSX1
XDFFPOSX1_130 MUX2X1_8/A NOR2X1_18/A NOR2X1_72/Y gnd vdd DFFPOSX1
XAND2X2_16 MUX2X1_6/B INVX1_48/A gnd OAI22X1_3/C vdd AND2X2
XCLKBUF1_14 reset gnd INVX2_11/A vdd CLKBUF1
XFILL_13_2_0 gnd vdd FILL
XNOR2X1_16 NOR2X1_18/A MUX2X1_5/Y gnd NOR2X1_16/Y vdd NOR2X1
XNOR2X1_38 NOR2X1_38/A NOR2X1_38/B gnd NOR2X1_38/Y vdd NOR2X1
XNOR2X1_27 NOR2X1_84/A NOR2X1_27/B gnd NOR2X1_27/Y vdd NOR2X1
XNOR2X1_49 INVX1_21/A INVX2_12/A gnd NOR2X1_49/Y vdd NOR2X1
XNAND3X1_16 INVX1_20/A INVX1_22/A NOR2X1_49/Y gnd OAI21X1_40/C vdd NAND3X1
XFILL_2_1_0 gnd vdd FILL
XMUX2X1_23 key[2] MUX2X1_3/A AND2X2_4/Y gnd NOR2X1_75/B vdd MUX2X1
XMUX2X1_45 MUX2X1_9/A MUX2X1_45/B BUFX4_3/Y gnd MUX2X1_45/Y vdd MUX2X1
XMUX2X1_34 MUX2X1_34/A MUX2X1_34/B BUFX4_3/Y gnd INVX1_39/A vdd MUX2X1
XFILL_10_0_0 gnd vdd FILL
XNOR2X1_106 NOR3X1_2/B NOR2X1_106/B gnd INVX1_5/A vdd NOR2X1
XMUX2X1_12 MUX2X1_46/A XOR2X1_7/A MUX2X1_9/S gnd NOR2X1_23/B vdd MUX2X1
XNAND2X1_60 INVX1_5/A NOR2X1_6/B gnd NOR2X1_107/B vdd NAND2X1
XINVX1_19 NOR3X1_5/Y gnd INVX1_19/Y vdd INVX1
XFILL_14_1 gnd vdd FILL
XFILL_7_0_0 gnd vdd FILL
XOAI21X1_25 BUFX4_10/Y MUX2X1_33/A INVX8_2/Y gnd OAI21X1_25/Y vdd OAI21X1
XOAI21X1_36 BUFX4_11/Y MUX2X1_7/A INVX8_2/Y gnd OAI21X1_36/Y vdd OAI21X1
XOAI21X1_47 INVX1_36/Y BUFX4_8/Y OAI21X1_47/C gnd OAI21X1_47/Y vdd OAI21X1
XOAI21X1_58 INVX1_49/Y BUFX4_8/Y OAI21X1_58/C gnd OAI21X1_58/Y vdd OAI21X1
XOAI21X1_14 OR2X2_2/A OR2X2_2/B INVX1_10/Y gnd NAND3X1_4/B vdd OAI21X1
XDFFPOSX1_142 MUX2X1_4/A CLKBUF1_1/Y NOR2X1_76/Y gnd vdd DFFPOSX1
XDFFPOSX1_120 MUX2X1_35/A NOR2X1_84/A NOR2X1_78/Y gnd vdd DFFPOSX1
XAND2X2_17 MUX2X1_9/B INVX2_2/A gnd OAI22X1_4/A vdd AND2X2
XDFFPOSX1_131 MUX2X1_9/A INVX8_2/A NOR2X1_81/Y gnd vdd DFFPOSX1
XCLKBUF1_15 reset gnd NOR2X1_75/A vdd CLKBUF1
XFILL_13_2_1 gnd vdd FILL
XXNOR2X1_1 OR2X2_2/A INVX2_2/Y gnd XNOR2X1_1/Y vdd XNOR2X1
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XAND2X2_1 OR2X2_1/Y AND2X2_1/B gnd AND2X2_1/Y vdd AND2X2
XFILL_2_1 gnd vdd FILL
XNOR2X1_28 INVX1_8/A INVX2_3/Y gnd NOR2X1_28/Y vdd NOR2X1
XNAND3X1_17 INVX2_10/A INVX1_20/A INVX1_21/A gnd XNOR2X1_6/A vdd NAND3X1
XNOR2X1_17 NOR2X1_25/A MUX2X1_6/Y gnd NOR2X1_17/Y vdd NOR2X1
XMUX2X1_24 key[3] MUX2X1_4/A AND2X2_4/Y gnd NOR2X1_76/B vdd MUX2X1
XMUX2X1_13 MUX2X1_33/A NOR2X1_86/A MUX2X1_9/S gnd NOR2X1_24/B vdd MUX2X1
XMUX2X1_35 MUX2X1_35/A MUX2X1_35/B BUFX4_3/Y gnd MUX2X1_35/Y vdd MUX2X1
XMUX2X1_46 MUX2X1_46/A MUX2X1_46/B BUFX4_1/Y gnd INVX1_57/A vdd MUX2X1
XFILL_10_0_1 gnd vdd FILL
XNOR2X1_39 INVX1_7/A INVX2_2/Y gnd NOR2X1_39/Y vdd NOR2X1
XNOR2X1_107 INVX2_15/Y NOR2X1_107/B gnd NOR2X1_107/Y vdd NOR2X1
XFILL_2_1_1 gnd vdd FILL
XNAND2X1_50 OAI21X1_2/B AOI21X1_4/C gnd NOR2X1_102/A vdd NAND2X1
XFILL_14_2 gnd vdd FILL
XOAI21X1_26 XNOR2X1_3/A INVX4_1/Y INVX1_12/Y gnd NAND3X1_7/C vdd OAI21X1
XOAI21X1_37 XNOR2X1_5/A INVX2_7/Y INVX1_16/Y gnd OAI21X1_37/Y vdd OAI21X1
XOAI21X1_59 INVX1_50/Y BUFX4_9/Y OAI21X1_59/C gnd OAI21X1_59/Y vdd OAI21X1
XOAI21X1_48 INVX1_37/Y BUFX4_8/Y OAI21X1_48/C gnd OAI21X1_48/Y vdd OAI21X1
XFILL_7_0_1 gnd vdd FILL
XOAI21X1_15 BUFX4_14/Y MUX2X1_48/A INVX8_2/Y gnd OAI21X1_15/Y vdd OAI21X1
XDFFPOSX1_143 MUX2X1_5/A CLKBUF1_1/Y NOR2X1_69/Y gnd vdd DFFPOSX1
XDFFPOSX1_121 MUX2X1_36/A NOR2X1_79/A NOR2X1_79/Y gnd vdd DFFPOSX1
XDFFPOSX1_132 MUX2X1_47/A NOR2X1_84/A NOR2X1_82/Y gnd vdd DFFPOSX1
XAND2X2_18 NOR2X1_99/A INVX1_7/A gnd OAI22X1_4/C vdd AND2X2
XDFFPOSX1_110 INVX1_24/A CLKBUF1_4/Y NOR2X1_60/Y gnd vdd DFFPOSX1
XCLKBUF1_16 reset gnd NOR2X1_79/A vdd CLKBUF1
XXNOR2X1_2 INVX1_41/A XNOR2X1_2/B gnd XNOR2X1_2/Y vdd XNOR2X1
XINVX1_2 INVX1_2/A gnd OR2X2_1/B vdd INVX1
XAND2X2_2 NOR3X1_2/Y AND2X2_2/B gnd AND2X2_2/Y vdd AND2X2
XNOR2X1_18 NOR2X1_18/A MUX2X1_7/Y gnd NOR2X1_18/Y vdd NOR2X1
XNOR2X1_29 INVX2_4/A INVX1_11/A gnd NOR2X1_29/Y vdd NOR2X1
XNAND3X1_18 INVX2_11/Y OAI21X1_40/C NOR3X1_6/Y gnd NOR2X1_53/B vdd NAND3X1
XMUX2X1_36 MUX2X1_36/A MUX2X1_36/B BUFX4_3/Y gnd NOR2X1_89/A vdd MUX2X1
XMUX2X1_25 MUX2X1_9/A MUX2X1_33/A AND2X2_4/Y gnd NOR2X1_77/B vdd MUX2X1
XMUX2X1_47 MUX2X1_47/A MUX2X1_47/B BUFX4_1/Y gnd MUX2X1_47/Y vdd MUX2X1
XMUX2X1_14 MUX2X1_35/A NOR2X1_87/A MUX2X1_9/S gnd NOR2X1_25/B vdd MUX2X1
XNAND2X1_40 XOR2X1_4/A BUFX4_6/Y gnd OAI21X1_53/C vdd NAND2X1
XNAND2X1_51 INVX1_1/A OAI21X1_4/B gnd NOR2X1_102/B vdd NAND2X1
XNOR2X1_108 OAI21X1_67/A INVX2_15/Y gnd NOR2X1_108/Y vdd NOR2X1
XOAI21X1_27 BUFX4_10/Y MUX2X1_35/A INVX8_2/Y gnd OAI21X1_27/Y vdd OAI21X1
XOAI21X1_49 INVX1_38/Y BUFX4_6/Y OAI21X1_49/C gnd OAI21X1_49/Y vdd OAI21X1
XOAI21X1_38 BUFX4_12/Y MUX2X1_8/A INVX8_2/Y gnd OAI21X1_38/Y vdd OAI21X1
XOAI21X1_16 OR2X2_2/Y NOR2X1_31/B BUFX4_14/Y gnd OAI21X1_16/Y vdd OAI21X1
XDFFPOSX1_144 MUX2X1_6/A CLKBUF1_3/Y NOR2X1_70/Y gnd vdd DFFPOSX1
XAND2X2_19 OAI21X1_2/B AOI21X1_4/C gnd AND2X2_19/Y vdd AND2X2
XDFFPOSX1_111 INVX2_13/A CLKBUF1_4/Y NOR2X1_61/Y gnd vdd DFFPOSX1
XDFFPOSX1_122 MUX2X1_34/A INVX8_2/A NOR2X1_80/Y gnd vdd DFFPOSX1
XDFFPOSX1_100 INVX1_22/A INVX2_11/A AOI21X1_26/Y gnd vdd DFFPOSX1
XDFFPOSX1_133 MUX2X1_48/A INVX8_2/A NOR2X1_83/Y gnd vdd DFFPOSX1
XFILL_0_2_0 gnd vdd FILL
XFILL_16_2_0 gnd vdd FILL
XCLKBUF1_17 reset gnd NOR2X1_77/A vdd CLKBUF1
XXNOR2X1_3 XNOR2X1_3/A INVX4_1/Y gnd XNOR2X1_3/Y vdd XNOR2X1
XOR2X2_1 OR2X2_1/A OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XFILL_13_0_0 gnd vdd FILL
XFILL_5_1_0 gnd vdd FILL
XAND2X2_3 key[1] key[3] gnd AND2X2_3/Y vdd AND2X2
XNAND3X1_19 INVX1_23/A INVX1_25/A NOR2X1_56/Y gnd OAI21X1_43/C vdd NAND3X1
XNOR2X1_19 NOR2X1_25/A MUX2X1_8/Y gnd NOR2X1_19/Y vdd NOR2X1
XMUX2X1_48 MUX2X1_48/A MUX2X1_48/B BUFX4_1/Y gnd MUX2X1_48/Y vdd MUX2X1
XMUX2X1_37 MUX2X1_1/A MUX2X1_37/B BUFX4_4/Y gnd NOR2X1_92/A vdd MUX2X1
XMUX2X1_26 MUX2X1_47/A MUX2X1_35/A AND2X2_4/Y gnd NOR2X1_78/B vdd MUX2X1
XMUX2X1_15 MUX2X1_36/A XOR2X1_2/A MUX2X1_9/S gnd NOR2X1_26/B vdd MUX2X1
XNOR2X1_109 INVX2_17/Y OAI21X1_67/Y gnd NOR2X1_109/Y vdd NOR2X1
XNAND2X1_41 XOR2X1_3/A BUFX4_6/Y gnd OAI21X1_54/C vdd NAND2X1
XNAND2X1_52 OAI21X1_67/A OAI21X1_67/B gnd OR2X2_10/A vdd NAND2X1
XNAND2X1_30 OAI21X1_40/C OAI21X1_43/C gnd INVX1_27/A vdd NAND2X1
XOAI22X1_1 OAI22X1_1/A OAI22X1_1/B OAI22X1_1/C OAI22X1_1/D gnd NOR3X1_9/C vdd OAI22X1
XOAI21X1_28 NAND3X1_7/A NOR2X1_38/Y INVX2_5/Y gnd OAI21X1_29/C vdd OAI21X1
XOAI21X1_39 INVX2_8/Y NOR3X1_7/B INVX1_19/Y gnd BUFX4_4/A vdd OAI21X1
XINVX2_10 INVX2_10/A gnd INVX2_10/Y vdd INVX2
XOAI21X1_17 BUFX4_14/Y MUX2X1_46/A INVX8_2/Y gnd NOR2X1_33/A vdd OAI21X1
XFILL_12_1 gnd vdd FILL
XDFFPOSX1_123 MUX2X1_1/A NOR2X1_77/A NOR2X1_73/Y gnd vdd DFFPOSX1
XDFFPOSX1_145 MUX2X1_7/A CLKBUF1_3/Y NOR2X1_71/Y gnd vdd DFFPOSX1
XDFFPOSX1_134 MUX2X1_46/A INVX8_2/A NOR2X1_84/Y gnd vdd DFFPOSX1
XFILL_0_2_1 gnd vdd FILL
XDFFPOSX1_101 INVX1_20/A CLKBUF1_4/Y NOR2X1_52/Y gnd vdd DFFPOSX1
XDFFPOSX1_112 INVX1_25/A CLKBUF1_5/Y AOI21X1_27/Y gnd vdd DFFPOSX1
XFILL_16_2_1 gnd vdd FILL
XXNOR2X1_4 XNOR2X1_4/A INVX2_6/Y gnd XNOR2X1_4/Y vdd XNOR2X1
XCLKBUF1_18 reset gnd NOR2X1_18/A vdd CLKBUF1
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XFILL_5_1_1 gnd vdd FILL
XFILL_13_0_1 gnd vdd FILL
XAND2X2_4 AND2X2_4/A OR2X2_9/A gnd AND2X2_4/Y vdd AND2X2
XMUX2X1_27 MUX2X1_48/A MUX2X1_36/A AND2X2_4/Y gnd NOR2X1_79/B vdd MUX2X1
XMUX2X1_38 MUX2X1_4/A MUX2X1_38/B BUFX4_4/Y gnd INVX1_45/A vdd MUX2X1
XMUX2X1_16 MUX2X1_34/A XOR2X1_1/A MUX2X1_9/S gnd NOR2X1_27/B vdd MUX2X1
XNAND2X1_20 NOR2X1_44/Y AND2X2_3/Y gnd INVX1_26/A vdd NAND2X1
XNAND2X1_42 MUX2X1_5/B BUFX4_9/Y gnd OAI21X1_56/C vdd NAND2X1
XNAND2X1_53 AOI21X1_2/C AOI21X1_2/A gnd OR2X2_10/B vdd NAND2X1
XNAND2X1_31 INVX2_14/Y INVX1_32/Y gnd NAND2X1_31/Y vdd NAND2X1
XOAI22X1_2 OAI22X1_2/A OAI22X1_2/B OAI22X1_2/C OAI22X1_2/D gnd OAI22X1_2/Y vdd OAI22X1
XINVX2_11 INVX2_11/A gnd INVX2_11/Y vdd INVX2
XOAI21X1_18 BUFX4_13/Y MUX2X1_1/A INVX8_2/Y gnd OAI21X1_18/Y vdd OAI21X1
XOAI21X1_29 INVX2_5/Y NAND3X1_7/A OAI21X1_29/C gnd OAI21X1_29/Y vdd OAI21X1
XDFFPOSX1_124 MUX2X1_2/A NOR2X1_75/A NOR2X1_74/Y gnd vdd DFFPOSX1
XDFFPOSX1_135 MUX2X1_33/A CLKBUF1_1/Y NOR2X1_77/Y gnd vdd DFFPOSX1
XDFFPOSX1_146 MUX2X1_8/A CLKBUF1_3/Y NOR2X1_72/Y gnd vdd DFFPOSX1
XFILL_12_2 gnd vdd FILL
XDFFPOSX1_102 INVX1_21/A CLKBUF1_2/Y NOR2X1_53/Y gnd vdd DFFPOSX1
XDFFPOSX1_113 NOR3X1_7/B NOR2X1_104/A AOI21X1_29/Y gnd vdd DFFPOSX1
XOR2X2_10 OR2X2_10/A OR2X2_10/B gnd OR2X2_10/Y vdd OR2X2
XXNOR2X1_5 XNOR2X1_5/A INVX2_7/Y gnd XNOR2X1_5/Y vdd XNOR2X1
XOR2X2_3 OR2X2_3/A OR2X2_3/B gnd OR2X2_3/Y vdd OR2X2
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
.ends

