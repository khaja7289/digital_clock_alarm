module alarm_clock_top (clock, key[0], key[1], key[2], key[3], reset, time_button, alarm_button, fastwatch, ms_hour[0], ms_hour[1], ms_hour[2], ms_hour[3], ms_hour[4], ms_hour[5], ms_hour[6], ms_hour[7], ls_hour[0], ls_hour[1], ls_hour[2], ls_hour[3], ls_hour[4], ls_hour[5], ls_hour[6], ls_hour[7], ms_minute[0], ms_minute[1], ms_minute[2], ms_minute[3], ms_minute[4], ms_minute[5], ms_minute[6], ms_minute[7], ls_minute[0], ls_minute[1], ls_minute[2], ls_minute[3], ls_minute[4], ls_minute[5], ls_minute[6], ls_minute[7], alarm_sound);

input clock;
input key[0];
input key[1];
input key[2];
input key[3];
input reset;
input time_button;
input alarm_button;
input fastwatch;
output ms_hour[0];
output ms_hour[1];
output ms_hour[2];
output ms_hour[3];
output ms_hour[4];
output ms_hour[5];
output ms_hour[6];
output ms_hour[7];
output ls_hour[0];
output ls_hour[1];
output ls_hour[2];
output ls_hour[3];
output ls_hour[4];
output ls_hour[5];
output ls_hour[6];
output ls_hour[7];
output ms_minute[0];
output ms_minute[1];
output ms_minute[2];
output ms_minute[3];
output ms_minute[4];
output ms_minute[5];
output ms_minute[6];
output ms_minute[7];
output ls_minute[0];
output ls_minute[1];
output ls_minute[2];
output ls_minute[3];
output ls_minute[4];
output ls_minute[5];
output ls_minute[6];
output ls_minute[7];
output alarm_sound;

BUFX4 BUFX4_1 ( .A(fsm1_show_new_time), .Y(fsm1_show_new_time_bF_buf3) );
BUFX4 BUFX4_2 ( .A(fsm1_show_new_time), .Y(fsm1_show_new_time_bF_buf2) );
BUFX4 BUFX4_3 ( .A(fsm1_show_new_time), .Y(fsm1_show_new_time_bF_buf1) );
BUFX4 BUFX4_4 ( .A(fsm1_show_new_time), .Y(fsm1_show_new_time_bF_buf0) );
CLKBUF1 CLKBUF1_1 ( .A(clock), .Y(clock_bF_buf7) );
CLKBUF1 CLKBUF1_2 ( .A(clock), .Y(clock_bF_buf6) );
CLKBUF1 CLKBUF1_3 ( .A(clock), .Y(clock_bF_buf5) );
CLKBUF1 CLKBUF1_4 ( .A(clock), .Y(clock_bF_buf4) );
CLKBUF1 CLKBUF1_5 ( .A(clock), .Y(clock_bF_buf3) );
CLKBUF1 CLKBUF1_6 ( .A(clock), .Y(clock_bF_buf2) );
CLKBUF1 CLKBUF1_7 ( .A(clock), .Y(clock_bF_buf1) );
CLKBUF1 CLKBUF1_8 ( .A(clock), .Y(clock_bF_buf0) );
BUFX4 BUFX4_5 ( .A(fsm1__25_), .Y(fsm1__25__bF_buf4) );
BUFX4 BUFX4_6 ( .A(fsm1__25_), .Y(fsm1__25__bF_buf3) );
BUFX4 BUFX4_7 ( .A(fsm1__25_), .Y(fsm1__25__bF_buf2) );
BUFX4 BUFX4_8 ( .A(fsm1__25_), .Y(fsm1__25__bF_buf1) );
BUFX4 BUFX4_9 ( .A(fsm1__25_), .Y(fsm1__25__bF_buf0) );
BUFX4 BUFX4_10 ( .A(_84_), .Y(_84__bF_buf4) );
BUFX4 BUFX4_11 ( .A(_84_), .Y(_84__bF_buf3) );
BUFX4 BUFX4_12 ( .A(_84_), .Y(_84__bF_buf2) );
BUFX4 BUFX4_13 ( .A(_84_), .Y(_84__bF_buf1) );
BUFX4 BUFX4_14 ( .A(_84_), .Y(_84__bF_buf0) );
CLKBUF1 CLKBUF1_9 ( .A(reset), .Y(reset_bF_buf9) );
CLKBUF1 CLKBUF1_10 ( .A(reset), .Y(reset_bF_buf8) );
CLKBUF1 CLKBUF1_11 ( .A(reset), .Y(reset_bF_buf7) );
CLKBUF1 CLKBUF1_12 ( .A(reset), .Y(reset_bF_buf6) );
CLKBUF1 CLKBUF1_13 ( .A(reset), .Y(reset_bF_buf5) );
CLKBUF1 CLKBUF1_14 ( .A(reset), .Y(reset_bF_buf4) );
CLKBUF1 CLKBUF1_15 ( .A(reset), .Y(reset_bF_buf3) );
CLKBUF1 CLKBUF1_16 ( .A(reset), .Y(reset_bF_buf2) );
CLKBUF1 CLKBUF1_17 ( .A(reset), .Y(reset_bF_buf1) );
CLKBUF1 CLKBUF1_18 ( .A(reset), .Y(reset_bF_buf0) );
AOI21X1 AOI21X1_1 ( .A(tgen1_count_2_), .B(_339_), .C(_341_), .Y(tgen1__00__2_) );
AOI21X1 AOI21X1_2 ( .A(tgen1_count_2_), .B(_339_), .C(tgen1_count_3_), .Y(_342_) );
OAI21X1 OAI21X1_1 ( .A(_320_), .B(_321_), .C(_324_), .Y(_343_) );
NOR2X1 NOR2X1_1 ( .A(_343_), .B(_342_), .Y(tgen1__00__3_) );
NAND2X1 NAND2X1_1 ( .A(tgen1_count_4_), .B(_322_), .Y(_344_) );
INVX2 INVX2_1 ( .A(_344_), .Y(_345_) );
OAI21X1 OAI21X1_2 ( .A(_322_), .B(tgen1_count_4_), .C(_324_), .Y(_346_) );
NOR2X1 NOR2X1_2 ( .A(_346_), .B(_345_), .Y(tgen1__00__4_) );
INVX1 INVX1_1 ( .A(tgen1_count_5_), .Y(_347_) );
NOR2X1 NOR2X1_3 ( .A(_347_), .B(_344_), .Y(_348_) );
OAI21X1 OAI21X1_3 ( .A(_345_), .B(tgen1_count_5_), .C(_324_), .Y(_349_) );
NOR2X1 NOR2X1_4 ( .A(_348_), .B(_349_), .Y(tgen1__00__5_) );
OAI21X1 OAI21X1_4 ( .A(_348_), .B(tgen1_count_6_), .C(_324_), .Y(_350_) );
AOI21X1 AOI21X1_3 ( .A(_329_), .B(_345_), .C(_350_), .Y(tgen1__00__6_) );
AOI21X1 AOI21X1_4 ( .A(_329_), .B(_345_), .C(tgen1_count_7_), .Y(_351_) );
OAI21X1 OAI21X1_5 ( .A(_331_), .B(_330_), .C(_324_), .Y(_352_) );
NOR2X1 NOR2X1_5 ( .A(_352_), .B(_351_), .Y(tgen1__00__7_) );
INVX1 INVX1_2 ( .A(tgen1_count_8_), .Y(_353_) );
OR2X2 OR2X2_1 ( .A(_323_), .B(_353_), .Y(_354_) );
AOI21X1 AOI21X1_5 ( .A(_353_), .B(_323_), .C(_325_), .Y(_355_) );
AND2X2 AND2X2_1 ( .A(_354_), .B(_355_), .Y(tgen1__00__8_) );
INVX1 INVX1_3 ( .A(tgen1_count_9_), .Y(_356_) );
OAI21X1 OAI21X1_6 ( .A(_323_), .B(_332_), .C(_324_), .Y(_357_) );
AOI21X1 AOI21X1_6 ( .A(_356_), .B(_354_), .C(_357_), .Y(tgen1__00__9_) );
NOR2X1 NOR2X1_6 ( .A(tgen1_count_10_), .B(_333_), .Y(_358_) );
INVX1 INVX1_4 ( .A(_332_), .Y(_359_) );
NAND3X1 NAND3X1_1 ( .A(_359_), .B(_319_), .C(_322_), .Y(_360_) );
NOR2X1 NOR2X1_7 ( .A(_335_), .B(_360_), .Y(_361_) );
INVX1 INVX1_5 ( .A(_337_), .Y(_362_) );
OAI21X1 OAI21X1_7 ( .A(_362_), .B(_360_), .C(_324_), .Y(_363_) );
NOR3X1 NOR3X1_1 ( .A(_363_), .B(_361_), .C(_358_), .Y(tgen1__00__10_) );
NOR2X1 NOR2X1_8 ( .A(tgen1_count_11_), .B(_361_), .Y(_364_) );
INVX1 INVX1_6 ( .A(tgen1_count_11_), .Y(_365_) );
NAND2X1 NAND2X1_2 ( .A(tgen1_count_10_), .B(_333_), .Y(_309_) );
AOI21X1 AOI21X1_7 ( .A(_337_), .B(_333_), .C(_325_), .Y(_310_) );
OAI21X1 OAI21X1_8 ( .A(_365_), .B(_309_), .C(_310_), .Y(_311_) );
NOR2X1 NOR2X1_9 ( .A(_364_), .B(_311_), .Y(tgen1__00__11_) );
AOI21X1 AOI21X1_8 ( .A(tgen1_count_11_), .B(_361_), .C(tgen1_count_12_), .Y(_312_) );
OAI21X1 OAI21X1_9 ( .A(_334_), .B(_309_), .C(_310_), .Y(_313_) );
NOR2X1 NOR2X1_10 ( .A(_312_), .B(_313_), .Y(tgen1__00__12_) );
NOR3X1 NOR3X1_2 ( .A(_335_), .B(_334_), .C(_360_), .Y(_314_) );
AND2X2 AND2X2_2 ( .A(_314_), .B(tgen1_count_13_), .Y(_315_) );
OAI21X1 OAI21X1_10 ( .A(tgen1_count_13_), .B(_314_), .C(_310_), .Y(_316_) );
NOR2X1 NOR2X1_11 ( .A(_315_), .B(_316_), .Y(tgen1__00__13_) );
DFFPOSX1 DFFPOSX1_1 ( .CLK(reset_bF_buf9), .D(tgen1__03_), .Q(fsm1_one_second) );
DFFPOSX1 DFFPOSX1_2 ( .CLK(clock_bF_buf7), .D(tgen1__03_), .Q(fsm1_one_second) );
DFFPOSX1 DFFPOSX1_3 ( .CLK(reset_bF_buf8), .D(tgen1__00__0_), .Q(tgen1_count_0_) );
DFFPOSX1 DFFPOSX1_4 ( .CLK(reset_bF_buf7), .D(tgen1__00__1_), .Q(tgen1_count_1_) );
DFFPOSX1 DFFPOSX1_5 ( .CLK(reset_bF_buf6), .D(tgen1__00__2_), .Q(tgen1_count_2_) );
DFFPOSX1 DFFPOSX1_6 ( .CLK(reset_bF_buf5), .D(tgen1__00__3_), .Q(tgen1_count_3_) );
DFFPOSX1 DFFPOSX1_7 ( .CLK(reset_bF_buf4), .D(tgen1__00__4_), .Q(tgen1_count_4_) );
DFFPOSX1 DFFPOSX1_8 ( .CLK(reset_bF_buf3), .D(tgen1__00__5_), .Q(tgen1_count_5_) );
DFFPOSX1 DFFPOSX1_9 ( .CLK(reset_bF_buf2), .D(tgen1__00__6_), .Q(tgen1_count_6_) );
DFFPOSX1 DFFPOSX1_10 ( .CLK(reset_bF_buf1), .D(tgen1__00__7_), .Q(tgen1_count_7_) );
DFFPOSX1 DFFPOSX1_11 ( .CLK(reset_bF_buf0), .D(tgen1__00__8_), .Q(tgen1_count_8_) );
DFFPOSX1 DFFPOSX1_12 ( .CLK(reset_bF_buf9), .D(tgen1__00__9_), .Q(tgen1_count_9_) );
DFFPOSX1 DFFPOSX1_13 ( .CLK(reset_bF_buf8), .D(tgen1__00__10_), .Q(tgen1_count_10_) );
DFFPOSX1 DFFPOSX1_14 ( .CLK(reset_bF_buf7), .D(tgen1__00__11_), .Q(tgen1_count_11_) );
DFFPOSX1 DFFPOSX1_15 ( .CLK(reset_bF_buf6), .D(tgen1__00__12_), .Q(tgen1_count_12_) );
DFFPOSX1 DFFPOSX1_16 ( .CLK(reset_bF_buf5), .D(tgen1__00__13_), .Q(tgen1_count_13_) );
DFFPOSX1 DFFPOSX1_17 ( .CLK(reset_bF_buf4), .D(tgen1__02_), .Q(tgen1_one_minute_reg) );
DFFPOSX1 DFFPOSX1_18 ( .CLK(clock_bF_buf6), .D(tgen1__00__0_), .Q(tgen1_count_0_) );
DFFPOSX1 DFFPOSX1_19 ( .CLK(clock_bF_buf5), .D(tgen1__00__1_), .Q(tgen1_count_1_) );
DFFPOSX1 DFFPOSX1_20 ( .CLK(clock_bF_buf4), .D(tgen1__00__2_), .Q(tgen1_count_2_) );
DFFPOSX1 DFFPOSX1_21 ( .CLK(clock_bF_buf3), .D(tgen1__00__3_), .Q(tgen1_count_3_) );
DFFPOSX1 DFFPOSX1_22 ( .CLK(clock_bF_buf2), .D(tgen1__00__4_), .Q(tgen1_count_4_) );
DFFPOSX1 DFFPOSX1_23 ( .CLK(clock_bF_buf1), .D(tgen1__00__5_), .Q(tgen1_count_5_) );
DFFPOSX1 DFFPOSX1_24 ( .CLK(clock_bF_buf0), .D(tgen1__00__6_), .Q(tgen1_count_6_) );
DFFPOSX1 DFFPOSX1_25 ( .CLK(clock_bF_buf7), .D(tgen1__00__7_), .Q(tgen1_count_7_) );
DFFPOSX1 DFFPOSX1_26 ( .CLK(clock_bF_buf6), .D(tgen1__00__8_), .Q(tgen1_count_8_) );
DFFPOSX1 DFFPOSX1_27 ( .CLK(clock_bF_buf5), .D(tgen1__00__9_), .Q(tgen1_count_9_) );
DFFPOSX1 DFFPOSX1_28 ( .CLK(clock_bF_buf4), .D(tgen1__00__10_), .Q(tgen1_count_10_) );
DFFPOSX1 DFFPOSX1_29 ( .CLK(clock_bF_buf3), .D(tgen1__00__11_), .Q(tgen1_count_11_) );
DFFPOSX1 DFFPOSX1_30 ( .CLK(clock_bF_buf2), .D(tgen1__00__12_), .Q(tgen1_count_12_) );
DFFPOSX1 DFFPOSX1_31 ( .CLK(clock_bF_buf1), .D(tgen1__00__13_), .Q(tgen1_count_13_) );
DFFPOSX1 DFFPOSX1_32 ( .CLK(clock_bF_buf0), .D(tgen1__02_), .Q(tgen1_one_minute_reg) );
BUFX2 BUFX2_1 ( .A(_0_), .Y(alarm_sound) );
BUFX2 BUFX2_2 ( .A(_1__0_), .Y(ls_hour[0]) );
BUFX2 BUFX2_3 ( .A(_1__1_), .Y(ls_hour[1]) );
BUFX2 BUFX2_4 ( .A(_1__2_), .Y(ls_hour[2]) );
BUFX2 BUFX2_5 ( .A(_1__3_), .Y(ls_hour[3]) );
BUFX2 BUFX2_6 ( .A(1'b1), .Y(ls_hour[4]) );
BUFX2 BUFX2_7 ( .A(1'b1), .Y(ls_hour[5]) );
BUFX2 BUFX2_8 ( .A(1'b0), .Y(ls_hour[6]) );
BUFX2 BUFX2_9 ( .A(1'b0), .Y(ls_hour[7]) );
BUFX2 BUFX2_10 ( .A(_2__0_), .Y(ls_minute[0]) );
BUFX2 BUFX2_11 ( .A(_2__1_), .Y(ls_minute[1]) );
BUFX2 BUFX2_12 ( .A(_2__2_), .Y(ls_minute[2]) );
BUFX2 BUFX2_13 ( .A(_2__3_), .Y(ls_minute[3]) );
BUFX2 BUFX2_14 ( .A(1'b1), .Y(ls_minute[4]) );
BUFX2 BUFX2_15 ( .A(1'b1), .Y(ls_minute[5]) );
BUFX2 BUFX2_16 ( .A(1'b0), .Y(ls_minute[6]) );
BUFX2 BUFX2_17 ( .A(1'b0), .Y(ls_minute[7]) );
BUFX2 BUFX2_18 ( .A(_3__0_), .Y(ms_hour[0]) );
BUFX2 BUFX2_19 ( .A(_3__1_), .Y(ms_hour[1]) );
BUFX2 BUFX2_20 ( .A(_3__2_), .Y(ms_hour[2]) );
BUFX2 BUFX2_21 ( .A(_3__3_), .Y(ms_hour[3]) );
BUFX2 BUFX2_22 ( .A(1'b1), .Y(ms_hour[4]) );
BUFX2 BUFX2_23 ( .A(1'b1), .Y(ms_hour[5]) );
BUFX2 BUFX2_24 ( .A(1'b0), .Y(ms_hour[6]) );
BUFX2 BUFX2_25 ( .A(1'b0), .Y(ms_hour[7]) );
BUFX2 BUFX2_26 ( .A(_4__0_), .Y(ms_minute[0]) );
BUFX2 BUFX2_27 ( .A(_4__1_), .Y(ms_minute[1]) );
BUFX2 BUFX2_28 ( .A(_4__2_), .Y(ms_minute[2]) );
BUFX2 BUFX2_29 ( .A(_4__3_), .Y(ms_minute[3]) );
BUFX2 BUFX2_30 ( .A(1'b1), .Y(ms_minute[4]) );
BUFX2 BUFX2_31 ( .A(1'b1), .Y(ms_minute[5]) );
BUFX2 BUFX2_32 ( .A(1'b0), .Y(ms_minute[6]) );
BUFX2 BUFX2_33 ( .A(1'b0), .Y(ms_minute[7]) );
MUX2X1 MUX2X1_1 ( .A(alreg1_new_alarm_ls_min_0_), .B(alarm_time_ls_min_0_), .S(alreg1_load_new_alarm), .Y(_5_) );
NOR2X1 NOR2X1_12 ( .A(reset_bF_buf3), .B(_5_), .Y(alreg1__1__0_) );
MUX2X1 MUX2X1_2 ( .A(alreg1_new_alarm_ls_min_1_), .B(alarm_time_ls_min_1_), .S(alreg1_load_new_alarm), .Y(_6_) );
NOR2X1 NOR2X1_13 ( .A(reset_bF_buf2), .B(_6_), .Y(alreg1__1__1_) );
MUX2X1 MUX2X1_3 ( .A(alreg1_new_alarm_ls_min_2_), .B(alarm_time_ls_min_2_), .S(alreg1_load_new_alarm), .Y(_7_) );
NOR2X1 NOR2X1_14 ( .A(reset_bF_buf1), .B(_7_), .Y(alreg1__1__2_) );
MUX2X1 MUX2X1_4 ( .A(alreg1_new_alarm_ls_min_3_), .B(alarm_time_ls_min_3_), .S(alreg1_load_new_alarm), .Y(_8_) );
NOR2X1 NOR2X1_15 ( .A(reset_bF_buf0), .B(_8_), .Y(alreg1__1__3_) );
MUX2X1 MUX2X1_5 ( .A(alreg1_new_alarm_ms_hr_0_), .B(alarm_time_ms_hr_0_), .S(alreg1_load_new_alarm), .Y(_9_) );
NOR2X1 NOR2X1_16 ( .A(reset_bF_buf9), .B(_9_), .Y(alreg1__2__0_) );
MUX2X1 MUX2X1_6 ( .A(alreg1_new_alarm_ms_hr_1_), .B(alarm_time_ms_hr_1_), .S(alreg1_load_new_alarm), .Y(_10_) );
NOR2X1 NOR2X1_17 ( .A(reset_bF_buf8), .B(_10_), .Y(alreg1__2__1_) );
MUX2X1 MUX2X1_7 ( .A(alreg1_new_alarm_ms_hr_2_), .B(alarm_time_ms_hr_2_), .S(alreg1_load_new_alarm), .Y(_11_) );
NOR2X1 NOR2X1_18 ( .A(reset_bF_buf7), .B(_11_), .Y(alreg1__2__2_) );
MUX2X1 MUX2X1_8 ( .A(alreg1_new_alarm_ms_hr_3_), .B(alarm_time_ms_hr_3_), .S(alreg1_load_new_alarm), .Y(_12_) );
NOR2X1 NOR2X1_19 ( .A(reset_bF_buf6), .B(_12_), .Y(alreg1__2__3_) );
MUX2X1 MUX2X1_9 ( .A(alreg1_new_alarm_ms_min_0_), .B(alarm_time_ms_min_0_), .S(alreg1_load_new_alarm), .Y(_13_) );
NOR2X1 NOR2X1_20 ( .A(reset_bF_buf5), .B(_13_), .Y(alreg1__3__0_) );
MUX2X1 MUX2X1_10 ( .A(alreg1_new_alarm_ms_min_1_), .B(alarm_time_ms_min_1_), .S(alreg1_load_new_alarm), .Y(_14_) );
NOR2X1 NOR2X1_21 ( .A(reset_bF_buf4), .B(_14_), .Y(alreg1__3__1_) );
MUX2X1 MUX2X1_11 ( .A(alreg1_new_alarm_ms_min_2_), .B(alarm_time_ms_min_2_), .S(alreg1_load_new_alarm), .Y(_15_) );
NOR2X1 NOR2X1_22 ( .A(reset_bF_buf3), .B(_15_), .Y(alreg1__3__2_) );
MUX2X1 MUX2X1_12 ( .A(alreg1_new_alarm_ms_min_3_), .B(alarm_time_ms_min_3_), .S(alreg1_load_new_alarm), .Y(_16_) );
NOR2X1 NOR2X1_23 ( .A(reset_bF_buf2), .B(_16_), .Y(alreg1__3__3_) );
MUX2X1 MUX2X1_13 ( .A(alreg1_new_alarm_ls_hr_0_), .B(alarm_time_ls_hr_0_), .S(alreg1_load_new_alarm), .Y(_17_) );
NOR2X1 NOR2X1_24 ( .A(reset_bF_buf1), .B(_17_), .Y(alreg1__0__0_) );
MUX2X1 MUX2X1_14 ( .A(alreg1_new_alarm_ls_hr_1_), .B(alarm_time_ls_hr_1_), .S(alreg1_load_new_alarm), .Y(_18_) );
NOR2X1 NOR2X1_25 ( .A(reset_bF_buf0), .B(_18_), .Y(alreg1__0__1_) );
MUX2X1 MUX2X1_15 ( .A(alreg1_new_alarm_ls_hr_2_), .B(alarm_time_ls_hr_2_), .S(alreg1_load_new_alarm), .Y(_19_) );
NOR2X1 NOR2X1_26 ( .A(reset_bF_buf9), .B(_19_), .Y(alreg1__0__2_) );
MUX2X1 MUX2X1_16 ( .A(alreg1_new_alarm_ls_hr_3_), .B(alarm_time_ls_hr_3_), .S(alreg1_load_new_alarm), .Y(_20_) );
NOR2X1 NOR2X1_27 ( .A(reset_bF_buf8), .B(_20_), .Y(alreg1__0__3_) );
DFFPOSX1 DFFPOSX1_33 ( .CLK(reset_bF_buf7), .D(alreg1__3__0_), .Q(alarm_time_ms_min_0_) );
DFFPOSX1 DFFPOSX1_34 ( .CLK(reset_bF_buf6), .D(alreg1__3__1_), .Q(alarm_time_ms_min_1_) );
DFFPOSX1 DFFPOSX1_35 ( .CLK(reset_bF_buf5), .D(alreg1__3__2_), .Q(alarm_time_ms_min_2_) );
DFFPOSX1 DFFPOSX1_36 ( .CLK(reset_bF_buf4), .D(alreg1__3__3_), .Q(alarm_time_ms_min_3_) );
DFFPOSX1 DFFPOSX1_37 ( .CLK(reset_bF_buf3), .D(alreg1__0__0_), .Q(alarm_time_ls_hr_0_) );
DFFPOSX1 DFFPOSX1_38 ( .CLK(reset_bF_buf2), .D(alreg1__0__1_), .Q(alarm_time_ls_hr_1_) );
DFFPOSX1 DFFPOSX1_39 ( .CLK(reset_bF_buf1), .D(alreg1__0__2_), .Q(alarm_time_ls_hr_2_) );
DFFPOSX1 DFFPOSX1_40 ( .CLK(reset_bF_buf0), .D(alreg1__0__3_), .Q(alarm_time_ls_hr_3_) );
DFFPOSX1 DFFPOSX1_41 ( .CLK(reset_bF_buf9), .D(alreg1__1__0_), .Q(alarm_time_ls_min_0_) );
DFFPOSX1 DFFPOSX1_42 ( .CLK(reset_bF_buf8), .D(alreg1__1__1_), .Q(alarm_time_ls_min_1_) );
DFFPOSX1 DFFPOSX1_43 ( .CLK(reset_bF_buf7), .D(alreg1__1__2_), .Q(alarm_time_ls_min_2_) );
DFFPOSX1 DFFPOSX1_44 ( .CLK(reset_bF_buf6), .D(alreg1__1__3_), .Q(alarm_time_ls_min_3_) );
DFFPOSX1 DFFPOSX1_45 ( .CLK(reset_bF_buf5), .D(alreg1__2__0_), .Q(alarm_time_ms_hr_0_) );
DFFPOSX1 DFFPOSX1_46 ( .CLK(reset_bF_buf4), .D(alreg1__2__1_), .Q(alarm_time_ms_hr_1_) );
DFFPOSX1 DFFPOSX1_47 ( .CLK(reset_bF_buf3), .D(alreg1__2__2_), .Q(alarm_time_ms_hr_2_) );
DFFPOSX1 DFFPOSX1_48 ( .CLK(reset_bF_buf2), .D(alreg1__2__3_), .Q(alarm_time_ms_hr_3_) );
DFFPOSX1 DFFPOSX1_49 ( .CLK(clock_bF_buf7), .D(alreg1__3__0_), .Q(alarm_time_ms_min_0_) );
DFFPOSX1 DFFPOSX1_50 ( .CLK(clock_bF_buf6), .D(alreg1__3__1_), .Q(alarm_time_ms_min_1_) );
DFFPOSX1 DFFPOSX1_51 ( .CLK(clock_bF_buf5), .D(alreg1__3__2_), .Q(alarm_time_ms_min_2_) );
DFFPOSX1 DFFPOSX1_52 ( .CLK(clock_bF_buf4), .D(alreg1__3__3_), .Q(alarm_time_ms_min_3_) );
DFFPOSX1 DFFPOSX1_53 ( .CLK(clock_bF_buf3), .D(alreg1__0__0_), .Q(alarm_time_ls_hr_0_) );
DFFPOSX1 DFFPOSX1_54 ( .CLK(clock_bF_buf2), .D(alreg1__0__1_), .Q(alarm_time_ls_hr_1_) );
DFFPOSX1 DFFPOSX1_55 ( .CLK(clock_bF_buf1), .D(alreg1__0__2_), .Q(alarm_time_ls_hr_2_) );
DFFPOSX1 DFFPOSX1_56 ( .CLK(clock_bF_buf0), .D(alreg1__0__3_), .Q(alarm_time_ls_hr_3_) );
DFFPOSX1 DFFPOSX1_57 ( .CLK(clock_bF_buf7), .D(alreg1__1__0_), .Q(alarm_time_ls_min_0_) );
DFFPOSX1 DFFPOSX1_58 ( .CLK(clock_bF_buf6), .D(alreg1__1__1_), .Q(alarm_time_ls_min_1_) );
DFFPOSX1 DFFPOSX1_59 ( .CLK(clock_bF_buf5), .D(alreg1__1__2_), .Q(alarm_time_ls_min_2_) );
DFFPOSX1 DFFPOSX1_60 ( .CLK(clock_bF_buf4), .D(alreg1__1__3_), .Q(alarm_time_ls_min_3_) );
DFFPOSX1 DFFPOSX1_61 ( .CLK(clock_bF_buf3), .D(alreg1__2__0_), .Q(alarm_time_ms_hr_0_) );
DFFPOSX1 DFFPOSX1_62 ( .CLK(clock_bF_buf2), .D(alreg1__2__1_), .Q(alarm_time_ms_hr_1_) );
DFFPOSX1 DFFPOSX1_63 ( .CLK(clock_bF_buf1), .D(alreg1__2__2_), .Q(alarm_time_ms_hr_2_) );
DFFPOSX1 DFFPOSX1_64 ( .CLK(clock_bF_buf0), .D(alreg1__2__3_), .Q(alarm_time_ms_hr_3_) );
INVX8 INVX8_1 ( .A(count1_load_new_c), .Y(_84_) );
INVX2 INVX2_2 ( .A(count1_current_time_ms_min_0_), .Y(_85_) );
INVX2 INVX2_3 ( .A(count1_current_time_ls_min_3_), .Y(_86_) );
NOR2X1 NOR2X1_28 ( .A(count1_current_time_ls_min_2_), .B(_86_), .Y(_87_) );
NAND2X1 NAND2X1_3 ( .A(count1_current_time_ls_min_0_), .B(count1_one_minute), .Y(_88_) );
NOR2X1 NOR2X1_29 ( .A(count1_current_time_ls_min_1_), .B(_88_), .Y(_89_) );
NAND2X1 NAND2X1_4 ( .A(_87_), .B(_89_), .Y(_90_) );
XNOR2X1 XNOR2X1_1 ( .A(_90_), .B(_85_), .Y(_91_) );
INVX8 INVX8_2 ( .A(reset_bF_buf1), .Y(_92_) );
OAI21X1 OAI21X1_11 ( .A(_84__bF_buf4), .B(alreg1_new_alarm_ms_min_0_), .C(_92_), .Y(_93_) );
AOI21X1 AOI21X1_9 ( .A(_84__bF_buf3), .B(_91_), .C(_93_), .Y(count1__03__0_) );
INVX1 INVX1_7 ( .A(count1_current_time_ms_min_1_), .Y(_94_) );
OAI21X1 OAI21X1_12 ( .A(_90_), .B(_85_), .C(_94_), .Y(_95_) );
NAND2X1 NAND2X1_5 ( .A(count1_current_time_ms_min_0_), .B(count1_current_time_ms_min_1_), .Y(_96_) );
OR2X2 OR2X2_2 ( .A(_90_), .B(_96_), .Y(_97_) );
INVX1 INVX1_8 ( .A(count1_current_time_ls_min_2_), .Y(_98_) );
NAND2X1 NAND2X1_6 ( .A(count1_current_time_ls_min_3_), .B(_98_), .Y(_99_) );
INVX2 INVX2_4 ( .A(count1_current_time_ls_min_1_), .Y(_100_) );
NAND3X1 NAND3X1_2 ( .A(count1_current_time_ls_min_0_), .B(count1_one_minute), .C(_100_), .Y(_101_) );
NOR2X1 NOR2X1_30 ( .A(_99_), .B(_101_), .Y(_102_) );
NAND2X1 NAND2X1_7 ( .A(count1_current_time_ms_min_0_), .B(_94_), .Y(_103_) );
INVX1 INVX1_9 ( .A(count1_current_time_ms_min_3_), .Y(_104_) );
NAND2X1 NAND2X1_8 ( .A(count1_current_time_ms_min_2_), .B(_104_), .Y(_105_) );
NOR2X1 NOR2X1_31 ( .A(_103_), .B(_105_), .Y(_106_) );
NAND2X1 NAND2X1_9 ( .A(_106_), .B(_102_), .Y(_107_) );
NAND3X1 NAND3X1_3 ( .A(_95_), .B(_107_), .C(_97_), .Y(_108_) );
OAI21X1 OAI21X1_13 ( .A(_84__bF_buf2), .B(alreg1_new_alarm_ms_min_1_), .C(_92_), .Y(_109_) );
AOI21X1 AOI21X1_10 ( .A(_84__bF_buf1), .B(_108_), .C(_109_), .Y(count1__03__1_) );
NOR2X1 NOR2X1_32 ( .A(_96_), .B(_90_), .Y(_110_) );
NAND2X1 NAND2X1_10 ( .A(count1_current_time_ms_min_2_), .B(_110_), .Y(_111_) );
INVX1 INVX1_10 ( .A(count1_current_time_ms_min_2_), .Y(_112_) );
OAI21X1 OAI21X1_14 ( .A(_90_), .B(_96_), .C(_112_), .Y(_113_) );
NAND3X1 NAND3X1_4 ( .A(_107_), .B(_113_), .C(_111_), .Y(_114_) );
OAI21X1 OAI21X1_15 ( .A(_84__bF_buf0), .B(alreg1_new_alarm_ms_min_2_), .C(_92_), .Y(_115_) );
AOI21X1 AOI21X1_11 ( .A(_84__bF_buf4), .B(_114_), .C(_115_), .Y(count1__03__2_) );
OAI21X1 OAI21X1_16 ( .A(_97_), .B(_105_), .C(_84__bF_buf3), .Y(_116_) );
AOI21X1 AOI21X1_12 ( .A(count1_current_time_ms_min_3_), .B(_111_), .C(_116_), .Y(_117_) );
OAI21X1 OAI21X1_17 ( .A(_84__bF_buf2), .B(alreg1_new_alarm_ms_min_3_), .C(_92_), .Y(_118_) );
NOR2X1 NOR2X1_33 ( .A(_118_), .B(_117_), .Y(count1__03__3_) );
XNOR2X1 XNOR2X1_2 ( .A(count1_current_time_ls_min_0_), .B(count1_one_minute), .Y(_119_) );
OAI21X1 OAI21X1_18 ( .A(_84__bF_buf1), .B(alreg1_new_alarm_ls_min_0_), .C(_92_), .Y(_120_) );
AOI21X1 AOI21X1_13 ( .A(_84__bF_buf0), .B(_119_), .C(_120_), .Y(count1__01__0_) );
INVX1 INVX1_11 ( .A(_88_), .Y(_121_) );
OAI21X1 OAI21X1_19 ( .A(_121_), .B(_100_), .C(_84__bF_buf4), .Y(_122_) );
AOI21X1 AOI21X1_14 ( .A(_99_), .B(_89_), .C(_122_), .Y(_123_) );
OAI21X1 OAI21X1_20 ( .A(_84__bF_buf3), .B(alreg1_new_alarm_ls_min_1_), .C(_92_), .Y(_124_) );
NOR2X1 NOR2X1_34 ( .A(_124_), .B(_123_), .Y(count1__01__1_) );
NAND2X1 NAND2X1_11 ( .A(count1_current_time_ls_min_1_), .B(_121_), .Y(_125_) );
OR2X2 OR2X2_3 ( .A(_125_), .B(_98_), .Y(_21_) );
OAI21X1 OAI21X1_21 ( .A(_88_), .B(_100_), .C(_98_), .Y(_22_) );
NAND2X1 NAND2X1_12 ( .A(_22_), .B(_21_), .Y(_23_) );
OAI21X1 OAI21X1_22 ( .A(_84__bF_buf2), .B(alreg1_new_alarm_ls_min_2_), .C(_92_), .Y(_24_) );
AOI21X1 AOI21X1_15 ( .A(_84__bF_buf1), .B(_23_), .C(_24_), .Y(count1__01__2_) );
AOI21X1 AOI21X1_16 ( .A(_86_), .B(_21_), .C(_102_), .Y(_25_) );
OAI21X1 OAI21X1_23 ( .A(_86_), .B(_21_), .C(_25_), .Y(_26_) );
OAI21X1 OAI21X1_24 ( .A(_84__bF_buf0), .B(alreg1_new_alarm_ls_min_3_), .C(_92_), .Y(_27_) );
AOI21X1 AOI21X1_17 ( .A(_84__bF_buf4), .B(_26_), .C(_27_), .Y(count1__01__3_) );
INVX4 INVX4_1 ( .A(count1_current_time_ls_hr_0_), .Y(_28_) );
XNOR2X1 XNOR2X1_3 ( .A(_107_), .B(_28_), .Y(_29_) );
OAI21X1 OAI21X1_25 ( .A(_84__bF_buf3), .B(alreg1_new_alarm_ls_hr_0_), .C(_92_), .Y(_30_) );
AOI21X1 AOI21X1_18 ( .A(_84__bF_buf2), .B(_29_), .C(_30_), .Y(count1__00__0_) );
INVX1 INVX1_12 ( .A(count1_current_time_ls_hr_1_), .Y(_31_) );
OAI21X1 OAI21X1_26 ( .A(_107_), .B(_28_), .C(_31_), .Y(_32_) );
NOR2X1 NOR2X1_35 ( .A(_28_), .B(_31_), .Y(_33_) );
NAND3X1 NAND3X1_5 ( .A(_106_), .B(_33_), .C(_102_), .Y(_34_) );
NAND2X1 NAND2X1_13 ( .A(count1_current_time_ls_hr_0_), .B(_31_), .Y(_35_) );
INVX2 INVX2_5 ( .A(count1_current_time_ls_hr_2_), .Y(_36_) );
NAND2X1 NAND2X1_14 ( .A(count1_current_time_ls_hr_3_), .B(_36_), .Y(_37_) );
NOR2X1 NOR2X1_36 ( .A(_35_), .B(_37_), .Y(_38_) );
NAND3X1 NAND3X1_6 ( .A(_106_), .B(_38_), .C(_102_), .Y(_39_) );
NAND3X1 NAND3X1_7 ( .A(_34_), .B(_39_), .C(_32_), .Y(_40_) );
OAI21X1 OAI21X1_27 ( .A(_84__bF_buf1), .B(alreg1_new_alarm_ls_hr_1_), .C(_92_), .Y(_41_) );
AOI21X1 AOI21X1_19 ( .A(_84__bF_buf0), .B(_40_), .C(_41_), .Y(count1__00__1_) );
INVX1 INVX1_13 ( .A(count1_current_time_ls_hr_3_), .Y(_42_) );
NAND2X1 NAND2X1_15 ( .A(_36_), .B(_42_), .Y(_43_) );
INVX2 INVX2_6 ( .A(count1_current_time_ms_hr_0_), .Y(_44_) );
NOR2X1 NOR2X1_37 ( .A(count1_current_time_ms_hr_3_), .B(count1_current_time_ms_hr_2_), .Y(_45_) );
NAND3X1 NAND3X1_8 ( .A(_44_), .B(count1_current_time_ms_hr_1_), .C(_45_), .Y(_46_) );
NOR2X1 NOR2X1_38 ( .A(_43_), .B(_46_), .Y(_47_) );
OAI21X1 OAI21X1_28 ( .A(_34_), .B(_47_), .C(_36_), .Y(_48_) );
OAI21X1 OAI21X1_29 ( .A(_36_), .B(_34_), .C(_48_), .Y(_49_) );
OAI21X1 OAI21X1_30 ( .A(_84__bF_buf4), .B(alreg1_new_alarm_ls_hr_2_), .C(_92_), .Y(_50_) );
AOI21X1 AOI21X1_20 ( .A(_84__bF_buf3), .B(_49_), .C(_50_), .Y(count1__00__2_) );
NAND2X1 NAND2X1_16 ( .A(count1_current_time_ls_hr_2_), .B(_33_), .Y(_51_) );
OAI21X1 OAI21X1_31 ( .A(_107_), .B(_51_), .C(_42_), .Y(_52_) );
NOR2X1 NOR2X1_39 ( .A(count1_current_time_ms_min_1_), .B(_85_), .Y(_53_) );
NOR2X1 NOR2X1_40 ( .A(count1_current_time_ms_min_3_), .B(_112_), .Y(_54_) );
NAND2X1 NAND2X1_17 ( .A(_53_), .B(_54_), .Y(_55_) );
NOR2X1 NOR2X1_41 ( .A(_55_), .B(_90_), .Y(_56_) );
INVX1 INVX1_14 ( .A(_51_), .Y(_57_) );
NAND3X1 NAND3X1_9 ( .A(count1_current_time_ls_hr_3_), .B(_57_), .C(_56_), .Y(_58_) );
NAND3X1 NAND3X1_10 ( .A(_39_), .B(_52_), .C(_58_), .Y(_59_) );
OAI21X1 OAI21X1_32 ( .A(_84__bF_buf2), .B(alreg1_new_alarm_ls_hr_3_), .C(_92_), .Y(_60_) );
AOI21X1 AOI21X1_21 ( .A(_84__bF_buf1), .B(_59_), .C(_60_), .Y(count1__00__3_) );
XNOR2X1 XNOR2X1_4 ( .A(_39_), .B(_44_), .Y(_61_) );
OAI21X1 OAI21X1_33 ( .A(_84__bF_buf0), .B(alreg1_new_alarm_ms_hr_0_), .C(_92_), .Y(_62_) );
AOI21X1 AOI21X1_22 ( .A(_84__bF_buf4), .B(_61_), .C(_62_), .Y(count1__02__0_) );
INVX1 INVX1_15 ( .A(count1_current_time_ms_hr_1_), .Y(_63_) );
OAI21X1 OAI21X1_34 ( .A(_39_), .B(_44_), .C(_63_), .Y(_64_) );
NAND2X1 NAND2X1_18 ( .A(count1_current_time_ms_hr_0_), .B(count1_current_time_ms_hr_1_), .Y(_65_) );
NOR3X1 NOR3X1_3 ( .A(_35_), .B(_65_), .C(_37_), .Y(_66_) );
NAND3X1 NAND3X1_11 ( .A(_102_), .B(_106_), .C(_66_), .Y(_67_) );
NAND3X1 NAND3X1_12 ( .A(_33_), .B(_47_), .C(_56_), .Y(_68_) );
NAND3X1 NAND3X1_13 ( .A(_67_), .B(_68_), .C(_64_), .Y(_69_) );
OAI21X1 OAI21X1_35 ( .A(_84__bF_buf3), .B(alreg1_new_alarm_ms_hr_1_), .C(_92_), .Y(_70_) );
AOI21X1 AOI21X1_23 ( .A(_84__bF_buf2), .B(_69_), .C(_70_), .Y(count1__02__1_) );
INVX2 INVX2_7 ( .A(count1_current_time_ms_hr_2_), .Y(_71_) );
XNOR2X1 XNOR2X1_5 ( .A(_67_), .B(_71_), .Y(_72_) );
OAI21X1 OAI21X1_36 ( .A(_84__bF_buf1), .B(alreg1_new_alarm_ms_hr_2_), .C(_92_), .Y(_73_) );
AOI21X1 AOI21X1_24 ( .A(_84__bF_buf0), .B(_72_), .C(_73_), .Y(count1__02__2_) );
INVX1 INVX1_16 ( .A(count1_current_time_ms_hr_3_), .Y(_74_) );
OAI21X1 OAI21X1_37 ( .A(_67_), .B(_71_), .C(_74_), .Y(_75_) );
NOR2X1 NOR2X1_42 ( .A(count1_current_time_ls_hr_1_), .B(_28_), .Y(_76_) );
NOR2X1 NOR2X1_43 ( .A(count1_current_time_ls_hr_2_), .B(_42_), .Y(_77_) );
INVX1 INVX1_17 ( .A(_65_), .Y(_78_) );
NAND3X1 NAND3X1_14 ( .A(_78_), .B(_76_), .C(_77_), .Y(_79_) );
NOR3X1 NOR3X1_4 ( .A(_90_), .B(_55_), .C(_79_), .Y(_80_) );
NAND3X1 NAND3X1_15 ( .A(count1_current_time_ms_hr_3_), .B(count1_current_time_ms_hr_2_), .C(_80_), .Y(_81_) );
NAND2X1 NAND2X1_19 ( .A(_75_), .B(_81_), .Y(_82_) );
OAI21X1 OAI21X1_38 ( .A(_84__bF_buf4), .B(alreg1_new_alarm_ms_hr_3_), .C(_92_), .Y(_83_) );
AOI21X1 AOI21X1_25 ( .A(_84__bF_buf3), .B(_82_), .C(_83_), .Y(count1__02__3_) );
DFFPOSX1 DFFPOSX1_65 ( .CLK(reset_bF_buf0), .D(count1__00__0_), .Q(count1_current_time_ls_hr_0_) );
DFFPOSX1 DFFPOSX1_66 ( .CLK(reset_bF_buf9), .D(count1__00__1_), .Q(count1_current_time_ls_hr_1_) );
DFFPOSX1 DFFPOSX1_67 ( .CLK(reset_bF_buf8), .D(count1__00__2_), .Q(count1_current_time_ls_hr_2_) );
DFFPOSX1 DFFPOSX1_68 ( .CLK(reset_bF_buf7), .D(count1__00__3_), .Q(count1_current_time_ls_hr_3_) );
DFFPOSX1 DFFPOSX1_69 ( .CLK(reset_bF_buf6), .D(count1__01__0_), .Q(count1_current_time_ls_min_0_) );
DFFPOSX1 DFFPOSX1_70 ( .CLK(reset_bF_buf5), .D(count1__01__1_), .Q(count1_current_time_ls_min_1_) );
DFFPOSX1 DFFPOSX1_71 ( .CLK(reset_bF_buf4), .D(count1__01__2_), .Q(count1_current_time_ls_min_2_) );
DFFPOSX1 DFFPOSX1_72 ( .CLK(reset_bF_buf3), .D(count1__01__3_), .Q(count1_current_time_ls_min_3_) );
DFFPOSX1 DFFPOSX1_73 ( .CLK(reset_bF_buf2), .D(count1__02__0_), .Q(count1_current_time_ms_hr_0_) );
DFFPOSX1 DFFPOSX1_74 ( .CLK(reset_bF_buf1), .D(count1__02__1_), .Q(count1_current_time_ms_hr_1_) );
DFFPOSX1 DFFPOSX1_75 ( .CLK(reset_bF_buf0), .D(count1__02__2_), .Q(count1_current_time_ms_hr_2_) );
DFFPOSX1 DFFPOSX1_76 ( .CLK(reset_bF_buf9), .D(count1__02__3_), .Q(count1_current_time_ms_hr_3_) );
DFFPOSX1 DFFPOSX1_77 ( .CLK(reset_bF_buf8), .D(count1__03__0_), .Q(count1_current_time_ms_min_0_) );
DFFPOSX1 DFFPOSX1_78 ( .CLK(reset_bF_buf7), .D(count1__03__1_), .Q(count1_current_time_ms_min_1_) );
DFFPOSX1 DFFPOSX1_79 ( .CLK(reset_bF_buf6), .D(count1__03__2_), .Q(count1_current_time_ms_min_2_) );
DFFPOSX1 DFFPOSX1_80 ( .CLK(reset_bF_buf5), .D(count1__03__3_), .Q(count1_current_time_ms_min_3_) );
DFFPOSX1 DFFPOSX1_81 ( .CLK(clock_bF_buf7), .D(count1__00__0_), .Q(count1_current_time_ls_hr_0_) );
DFFPOSX1 DFFPOSX1_82 ( .CLK(clock_bF_buf6), .D(count1__00__1_), .Q(count1_current_time_ls_hr_1_) );
DFFPOSX1 DFFPOSX1_83 ( .CLK(clock_bF_buf5), .D(count1__00__2_), .Q(count1_current_time_ls_hr_2_) );
DFFPOSX1 DFFPOSX1_84 ( .CLK(clock_bF_buf4), .D(count1__00__3_), .Q(count1_current_time_ls_hr_3_) );
DFFPOSX1 DFFPOSX1_85 ( .CLK(clock_bF_buf3), .D(count1__01__0_), .Q(count1_current_time_ls_min_0_) );
DFFPOSX1 DFFPOSX1_86 ( .CLK(clock_bF_buf2), .D(count1__01__1_), .Q(count1_current_time_ls_min_1_) );
DFFPOSX1 DFFPOSX1_87 ( .CLK(clock_bF_buf1), .D(count1__01__2_), .Q(count1_current_time_ls_min_2_) );
DFFPOSX1 DFFPOSX1_88 ( .CLK(clock_bF_buf0), .D(count1__01__3_), .Q(count1_current_time_ls_min_3_) );
DFFPOSX1 DFFPOSX1_89 ( .CLK(clock_bF_buf7), .D(count1__02__0_), .Q(count1_current_time_ms_hr_0_) );
DFFPOSX1 DFFPOSX1_90 ( .CLK(clock_bF_buf6), .D(count1__02__1_), .Q(count1_current_time_ms_hr_1_) );
DFFPOSX1 DFFPOSX1_91 ( .CLK(clock_bF_buf5), .D(count1__02__2_), .Q(count1_current_time_ms_hr_2_) );
DFFPOSX1 DFFPOSX1_92 ( .CLK(clock_bF_buf4), .D(count1__02__3_), .Q(count1_current_time_ms_hr_3_) );
DFFPOSX1 DFFPOSX1_93 ( .CLK(clock_bF_buf3), .D(count1__03__0_), .Q(count1_current_time_ms_min_0_) );
DFFPOSX1 DFFPOSX1_94 ( .CLK(clock_bF_buf2), .D(count1__03__1_), .Q(count1_current_time_ms_min_1_) );
DFFPOSX1 DFFPOSX1_95 ( .CLK(clock_bF_buf1), .D(count1__03__2_), .Q(count1_current_time_ms_min_2_) );
DFFPOSX1 DFFPOSX1_96 ( .CLK(clock_bF_buf0), .D(count1__03__3_), .Q(count1_current_time_ms_min_3_) );
NOR2X1 NOR2X1_44 ( .A(key[0]), .B(key[2]), .Y(_194_) );
AND2X2 AND2X2_3 ( .A(key[1]), .B(key[3]), .Y(_195_) );
NAND2X1 NAND2X1_20 ( .A(_194_), .B(_195_), .Y(fsm1__39_) );
NAND2X1 NAND2X1_21 ( .A(fsm1_pre_state_1_), .B(fsm1_pre_state_0_), .Y(_196_) );
NOR2X1 NOR2X1_45 ( .A(fsm1_pre_state_2_), .B(_196_), .Y(fsm1__25_) );
INVX1 INVX1_18 ( .A(fsm1_pre_state_0_), .Y(_197_) );
NOR3X1 NOR3X1_5 ( .A(fsm1_pre_state_1_), .B(fsm1_pre_state_2_), .C(_197_), .Y(fsm1__22_) );
INVX2 INVX2_8 ( .A(fsm1_pre_state_1_), .Y(_198_) );
INVX2 INVX2_9 ( .A(fsm1_pre_state_2_), .Y(_199_) );
NOR3X1 NOR3X1_6 ( .A(_198_), .B(fsm1_pre_state_0_), .C(_199_), .Y(fsm1__24_) );
NOR2X1 NOR2X1_46 ( .A(fsm1_pre_state_0_), .B(_198_), .Y(_200_) );
AND2X2 AND2X2_4 ( .A(_200_), .B(_199_), .Y(fsm1_shift) );
NOR3X1 NOR3X1_7 ( .A(fsm1_pre_state_1_), .B(fsm1_pre_state_0_), .C(fsm1_pre_state_2_), .Y(_134_) );
NAND2X1 NAND2X1_22 ( .A(_198_), .B(_197_), .Y(_201_) );
NOR2X1 NOR2X1_47 ( .A(_199_), .B(_201_), .Y(alreg1_load_new_alarm) );
NAND2X1 NAND2X1_23 ( .A(fsm1_pre_state_0_), .B(_198_), .Y(_202_) );
NOR2X1 NOR2X1_48 ( .A(_199_), .B(_202_), .Y(count1_load_new_c) );
INVX1 INVX1_19 ( .A(fsm1__22_), .Y(_138_) );
OAI21X1 OAI21X1_39 ( .A(_198_), .B(fsm1_pre_state_0_), .C(_138_), .Y(fsm1_show_new_time) );
NOR2X1 NOR2X1_49 ( .A(fsm1_count2_1_), .B(fsm1_count2_2_), .Y(_139_) );
NAND3X1 NAND3X1_16 ( .A(fsm1_count2_0_), .B(fsm1_count2_3_), .C(_139_), .Y(_140_) );
INVX1 INVX1_20 ( .A(fsm1_count2_0_), .Y(_141_) );
NOR2X1 NOR2X1_50 ( .A(fsm1_one_second), .B(_141_), .Y(_142_) );
INVX2 INVX2_10 ( .A(fsm1_one_second), .Y(_143_) );
NOR2X1 NOR2X1_51 ( .A(fsm1_count2_0_), .B(_143_), .Y(_144_) );
OAI21X1 OAI21X1_40 ( .A(_142_), .B(_144_), .C(_140_), .Y(_145_) );
INVX2 INVX2_11 ( .A(reset_bF_buf4), .Y(_146_) );
NAND2X1 NAND2X1_24 ( .A(_146_), .B(fsm1__24_), .Y(_147_) );
NOR2X1 NOR2X1_52 ( .A(_147_), .B(_145_), .Y(fsm1__01__0_) );
INVX1 INVX1_21 ( .A(fsm1_count2_1_), .Y(_148_) );
OAI21X1 OAI21X1_41 ( .A(_143_), .B(_141_), .C(_148_), .Y(_149_) );
NAND3X1 NAND3X1_17 ( .A(fsm1_one_second), .B(fsm1_count2_0_), .C(fsm1_count2_1_), .Y(_150_) );
NAND2X1 NAND2X1_25 ( .A(_150_), .B(_149_), .Y(_151_) );
NAND3X1 NAND3X1_18 ( .A(_146_), .B(_140_), .C(fsm1__24_), .Y(_152_) );
NOR2X1 NOR2X1_53 ( .A(_151_), .B(_152_), .Y(fsm1__01__1_) );
INVX2 INVX2_12 ( .A(fsm1_count2_2_), .Y(_153_) );
XNOR2X1 XNOR2X1_6 ( .A(_150_), .B(_153_), .Y(_154_) );
NOR2X1 NOR2X1_54 ( .A(_154_), .B(_147_), .Y(fsm1__01__2_) );
OAI21X1 OAI21X1_42 ( .A(_150_), .B(_153_), .C(fsm1_count2_3_), .Y(_155_) );
INVX1 INVX1_22 ( .A(fsm1_count2_3_), .Y(_156_) );
NOR2X1 NOR2X1_55 ( .A(_153_), .B(_150_), .Y(_157_) );
NAND2X1 NAND2X1_26 ( .A(_156_), .B(_157_), .Y(_158_) );
AOI21X1 AOI21X1_26 ( .A(_155_), .B(_158_), .C(_152_), .Y(fsm1__01__3_) );
NOR2X1 NOR2X1_56 ( .A(fsm1_count1_1_), .B(fsm1_count1_2_), .Y(_159_) );
NAND3X1 NAND3X1_19 ( .A(fsm1_count1_0_), .B(fsm1_count1_3_), .C(_159_), .Y(_160_) );
NOR2X1 NOR2X1_57 ( .A(fsm1_count1_0_), .B(_143_), .Y(_161_) );
INVX1 INVX1_23 ( .A(fsm1_count1_0_), .Y(_162_) );
NOR2X1 NOR2X1_58 ( .A(fsm1_one_second), .B(_162_), .Y(_163_) );
OAI21X1 OAI21X1_43 ( .A(_161_), .B(_163_), .C(_160_), .Y(_164_) );
NAND2X1 NAND2X1_27 ( .A(_146_), .B(fsm1__22_), .Y(_165_) );
NOR2X1 NOR2X1_59 ( .A(_165_), .B(_164_), .Y(fsm1__00__0_) );
INVX1 INVX1_24 ( .A(fsm1_count1_1_), .Y(_166_) );
OAI21X1 OAI21X1_44 ( .A(_143_), .B(_162_), .C(_166_), .Y(_167_) );
NAND3X1 NAND3X1_20 ( .A(fsm1_one_second), .B(fsm1_count1_0_), .C(fsm1_count1_1_), .Y(_168_) );
NAND2X1 NAND2X1_28 ( .A(_168_), .B(_167_), .Y(_169_) );
NAND3X1 NAND3X1_21 ( .A(_146_), .B(fsm1__22_), .C(_160_), .Y(_170_) );
NOR2X1 NOR2X1_60 ( .A(_169_), .B(_170_), .Y(fsm1__00__1_) );
INVX2 INVX2_13 ( .A(fsm1_count1_2_), .Y(_171_) );
XNOR2X1 XNOR2X1_7 ( .A(_168_), .B(_171_), .Y(_172_) );
NOR2X1 NOR2X1_61 ( .A(_165_), .B(_172_), .Y(fsm1__00__2_) );
OAI21X1 OAI21X1_45 ( .A(_168_), .B(_171_), .C(fsm1_count1_3_), .Y(_173_) );
INVX1 INVX1_25 ( .A(fsm1_count1_3_), .Y(_174_) );
NOR2X1 NOR2X1_62 ( .A(_171_), .B(_168_), .Y(_175_) );
NAND2X1 NAND2X1_29 ( .A(_174_), .B(_175_), .Y(_176_) );
AOI21X1 AOI21X1_27 ( .A(_173_), .B(_176_), .C(_170_), .Y(fsm1__00__3_) );
INVX1 INVX1_26 ( .A(fsm1__39_), .Y(fsm1__19_) );
NAND2X1 NAND2X1_30 ( .A(_140_), .B(_160_), .Y(_177_) );
INVX1 INVX1_27 ( .A(_177_), .Y(_128__2_) );
INVX1 INVX1_28 ( .A(fsm1__13__0_), .Y(_178_) );
NOR2X1 NOR2X1_63 ( .A(_178_), .B(_177_), .Y(_131__0_) );
INVX1 INVX1_29 ( .A(fsm1__13__1_), .Y(_179_) );
NOR2X1 NOR2X1_64 ( .A(_179_), .B(_177_), .Y(_131__1_) );
INVX1 INVX1_30 ( .A(fsm1__13__2_), .Y(_180_) );
NOR2X1 NOR2X1_65 ( .A(_180_), .B(_177_), .Y(_131__2_) );
OR2X2 OR2X2_4 ( .A(fsm1__12__0_), .B(time_button), .Y(_130__0_) );
INVX1 INVX1_31 ( .A(time_button), .Y(_181_) );
AND2X2 AND2X2_5 ( .A(_181_), .B(fsm1__12__1_), .Y(_130__1_) );
OR2X2 OR2X2_5 ( .A(time_button), .B(fsm1__12__2_), .Y(_130__2_) );
INVX2 INVX2_14 ( .A(alarm_button), .Y(_182_) );
AND2X2 AND2X2_6 ( .A(_182_), .B(fsm1__11__0_), .Y(_129__0_) );
AND2X2 AND2X2_7 ( .A(_182_), .B(fsm1__11__1_), .Y(_129__1_) );
OR2X2 OR2X2_6 ( .A(alarm_button), .B(fsm1__11__2_), .Y(_129__2_) );
OR2X2 OR2X2_7 ( .A(fsm1__19_), .B(fsm1__09__0_), .Y(_127__0_) );
AND2X2 AND2X2_8 ( .A(fsm1__39_), .B(fsm1__09__2_), .Y(_127__2_) );
INVX1 INVX1_32 ( .A(fsm1__07__2_), .Y(_183_) );
NAND2X1 NAND2X1_31 ( .A(_182_), .B(_183_), .Y(_126__0_) );
OR2X2 OR2X2_8 ( .A(alarm_button), .B(fsm1__07__1_), .Y(_126__1_) );
NOR2X1 NOR2X1_66 ( .A(alarm_button), .B(_183_), .Y(_126__2_) );
INVX1 INVX1_33 ( .A(fsm1__04__1_), .Y(_184_) );
NOR3X1 NOR3X1_8 ( .A(fsm1_pre_state_2_), .B(_184_), .C(_196_), .Y(_185_) );
AOI21X1 AOI21X1_28 ( .A(fsm1__08__0_), .B(fsm1__24_), .C(_185_), .Y(_186_) );
AOI22X1 AOI22X1_1 ( .A(fsm1__06__0_), .B(_134_), .C(fsm1__22_), .D(fsm1__10__0_), .Y(_187_) );
AOI21X1 AOI21X1_29 ( .A(_187_), .B(_186_), .C(reset_bF_buf3), .Y(fsm1__03__0_) );
AOI21X1 AOI21X1_30 ( .A(fsm1__10__1_), .B(fsm1__22_), .C(_185_), .Y(_188_) );
OR2X2 OR2X2_9 ( .A(_199_), .B(fsm1__08__2_), .Y(_189_) );
AOI22X1 AOI22X1_2 ( .A(fsm1__06__1_), .B(_134_), .C(_189_), .D(_200_), .Y(_190_) );
AOI21X1 AOI21X1_31 ( .A(_190_), .B(_188_), .C(reset_bF_buf2), .Y(fsm1__03__1_) );
AOI22X1 AOI22X1_3 ( .A(fsm1__25__bF_buf4), .B(fsm1__04__2_), .C(fsm1__22_), .D(fsm1__10__2_), .Y(_191_) );
AOI22X1 AOI22X1_4 ( .A(fsm1__06__2_), .B(_134_), .C(_189_), .D(_200_), .Y(_192_) );
AOI21X1 AOI21X1_32 ( .A(_192_), .B(_191_), .C(reset_bF_buf1), .Y(fsm1__03__2_) );
AND2X2 AND2X2_9 ( .A(_134_), .B(_182_), .Y(_135_) );
AND2X2 AND2X2_10 ( .A(fsm1__24_), .B(fsm1__39_), .Y(_136_) );
NOR2X1 NOR2X1_67 ( .A(alarm_button), .B(_138_), .Y(_137_) );
NAND3X1 NAND3X1_22 ( .A(_181_), .B(_182_), .C(fsm1__22_), .Y(_193_) );
INVX1 INVX1_34 ( .A(_193_), .Y(_132_) );
NOR2X1 NOR2X1_68 ( .A(_177_), .B(_193_), .Y(_133_) );
DFFPOSX1 DFFPOSX1_97 ( .CLK(reset_bF_buf0), .D(fsm1__01__0_), .Q(fsm1_count2_0_) );
DFFPOSX1 DFFPOSX1_98 ( .CLK(reset_bF_buf9), .D(fsm1__01__1_), .Q(fsm1_count2_1_) );
DFFPOSX1 DFFPOSX1_99 ( .CLK(reset_bF_buf8), .D(fsm1__01__2_), .Q(fsm1_count2_2_) );
DFFPOSX1 DFFPOSX1_100 ( .CLK(reset_bF_buf7), .D(fsm1__01__3_), .Q(fsm1_count2_3_) );
DFFPOSX1 DFFPOSX1_101 ( .CLK(clock_bF_buf7), .D(fsm1__01__0_), .Q(fsm1_count2_0_) );
DFFPOSX1 DFFPOSX1_102 ( .CLK(clock_bF_buf6), .D(fsm1__01__1_), .Q(fsm1_count2_1_) );
DFFPOSX1 DFFPOSX1_103 ( .CLK(clock_bF_buf5), .D(fsm1__01__2_), .Q(fsm1_count2_2_) );
DFFPOSX1 DFFPOSX1_104 ( .CLK(clock_bF_buf4), .D(fsm1__01__3_), .Q(fsm1_count2_3_) );
DFFPOSX1 DFFPOSX1_105 ( .CLK(reset_bF_buf6), .D(fsm1__00__0_), .Q(fsm1_count1_0_) );
DFFPOSX1 DFFPOSX1_106 ( .CLK(reset_bF_buf5), .D(fsm1__00__1_), .Q(fsm1_count1_1_) );
DFFPOSX1 DFFPOSX1_107 ( .CLK(reset_bF_buf4), .D(fsm1__00__2_), .Q(fsm1_count1_2_) );
DFFPOSX1 DFFPOSX1_108 ( .CLK(reset_bF_buf3), .D(fsm1__00__3_), .Q(fsm1_count1_3_) );
DFFPOSX1 DFFPOSX1_109 ( .CLK(clock_bF_buf3), .D(fsm1__00__0_), .Q(fsm1_count1_0_) );
DFFPOSX1 DFFPOSX1_110 ( .CLK(clock_bF_buf2), .D(fsm1__00__1_), .Q(fsm1_count1_1_) );
DFFPOSX1 DFFPOSX1_111 ( .CLK(clock_bF_buf1), .D(fsm1__00__2_), .Q(fsm1_count1_2_) );
DFFPOSX1 DFFPOSX1_112 ( .CLK(clock_bF_buf0), .D(fsm1__00__3_), .Q(fsm1_count1_3_) );
DFFPOSX1 DFFPOSX1_113 ( .CLK(reset_bF_buf2), .D(fsm1__03__0_), .Q(fsm1_pre_state_0_) );
DFFPOSX1 DFFPOSX1_114 ( .CLK(reset_bF_buf1), .D(fsm1__03__1_), .Q(fsm1_pre_state_1_) );
DFFPOSX1 DFFPOSX1_115 ( .CLK(reset_bF_buf0), .D(fsm1__03__2_), .Q(fsm1_pre_state_2_) );
DFFPOSX1 DFFPOSX1_116 ( .CLK(clock_bF_buf7), .D(fsm1__03__0_), .Q(fsm1_pre_state_0_) );
DFFPOSX1 DFFPOSX1_117 ( .CLK(clock_bF_buf6), .D(fsm1__03__1_), .Q(fsm1_pre_state_1_) );
DFFPOSX1 DFFPOSX1_118 ( .CLK(clock_bF_buf5), .D(fsm1__03__2_), .Q(fsm1_pre_state_2_) );
MUX2X1 MUX2X1_17 ( .A(alreg1_new_alarm_ls_hr_0_), .B(alreg1_new_alarm_ms_hr_0_), .S(fsm1_shift), .Y(_203_) );
NOR2X1 NOR2X1_69 ( .A(reset_bF_buf9), .B(_203_), .Y(keyreg1__2__0_) );
MUX2X1 MUX2X1_18 ( .A(alreg1_new_alarm_ls_hr_1_), .B(alreg1_new_alarm_ms_hr_1_), .S(fsm1_shift), .Y(_204_) );
NOR2X1 NOR2X1_70 ( .A(reset_bF_buf8), .B(_204_), .Y(keyreg1__2__1_) );
MUX2X1 MUX2X1_19 ( .A(alreg1_new_alarm_ls_hr_2_), .B(alreg1_new_alarm_ms_hr_2_), .S(fsm1_shift), .Y(_205_) );
NOR2X1 NOR2X1_71 ( .A(reset_bF_buf7), .B(_205_), .Y(keyreg1__2__2_) );
MUX2X1 MUX2X1_20 ( .A(alreg1_new_alarm_ls_hr_3_), .B(alreg1_new_alarm_ms_hr_3_), .S(fsm1_shift), .Y(_206_) );
NOR2X1 NOR2X1_72 ( .A(reset_bF_buf6), .B(_206_), .Y(keyreg1__2__3_) );
MUX2X1 MUX2X1_21 ( .A(key[0]), .B(alreg1_new_alarm_ls_min_0_), .S(fsm1_shift), .Y(_207_) );
NOR2X1 NOR2X1_73 ( .A(reset_bF_buf5), .B(_207_), .Y(keyreg1__1__0_) );
MUX2X1 MUX2X1_22 ( .A(key[1]), .B(alreg1_new_alarm_ls_min_1_), .S(fsm1_shift), .Y(_208_) );
NOR2X1 NOR2X1_74 ( .A(reset_bF_buf4), .B(_208_), .Y(keyreg1__1__1_) );
MUX2X1 MUX2X1_23 ( .A(key[2]), .B(alreg1_new_alarm_ls_min_2_), .S(fsm1_shift), .Y(_209_) );
NOR2X1 NOR2X1_75 ( .A(reset_bF_buf3), .B(_209_), .Y(keyreg1__1__2_) );
MUX2X1 MUX2X1_24 ( .A(key[3]), .B(alreg1_new_alarm_ls_min_3_), .S(fsm1_shift), .Y(_210_) );
NOR2X1 NOR2X1_76 ( .A(reset_bF_buf2), .B(_210_), .Y(keyreg1__1__3_) );
MUX2X1 MUX2X1_25 ( .A(alreg1_new_alarm_ms_min_0_), .B(alreg1_new_alarm_ls_hr_0_), .S(fsm1_shift), .Y(_211_) );
NOR2X1 NOR2X1_77 ( .A(reset_bF_buf1), .B(_211_), .Y(keyreg1__0__0_) );
MUX2X1 MUX2X1_26 ( .A(alreg1_new_alarm_ms_min_1_), .B(alreg1_new_alarm_ls_hr_1_), .S(fsm1_shift), .Y(_212_) );
NOR2X1 NOR2X1_78 ( .A(reset_bF_buf0), .B(_212_), .Y(keyreg1__0__1_) );
MUX2X1 MUX2X1_27 ( .A(alreg1_new_alarm_ms_min_2_), .B(alreg1_new_alarm_ls_hr_2_), .S(fsm1_shift), .Y(_213_) );
NOR2X1 NOR2X1_79 ( .A(reset_bF_buf9), .B(_213_), .Y(keyreg1__0__2_) );
MUX2X1 MUX2X1_28 ( .A(alreg1_new_alarm_ms_min_3_), .B(alreg1_new_alarm_ls_hr_3_), .S(fsm1_shift), .Y(_214_) );
NOR2X1 NOR2X1_80 ( .A(reset_bF_buf8), .B(_214_), .Y(keyreg1__0__3_) );
MUX2X1 MUX2X1_29 ( .A(alreg1_new_alarm_ls_min_0_), .B(alreg1_new_alarm_ms_min_0_), .S(fsm1_shift), .Y(_215_) );
NOR2X1 NOR2X1_81 ( .A(reset_bF_buf7), .B(_215_), .Y(keyreg1__3__0_) );
MUX2X1 MUX2X1_30 ( .A(alreg1_new_alarm_ls_min_1_), .B(alreg1_new_alarm_ms_min_1_), .S(fsm1_shift), .Y(_216_) );
NOR2X1 NOR2X1_82 ( .A(reset_bF_buf6), .B(_216_), .Y(keyreg1__3__1_) );
MUX2X1 MUX2X1_31 ( .A(alreg1_new_alarm_ls_min_2_), .B(alreg1_new_alarm_ms_min_2_), .S(fsm1_shift), .Y(_217_) );
NOR2X1 NOR2X1_83 ( .A(reset_bF_buf5), .B(_217_), .Y(keyreg1__3__2_) );
MUX2X1 MUX2X1_32 ( .A(alreg1_new_alarm_ls_min_3_), .B(alreg1_new_alarm_ms_min_3_), .S(fsm1_shift), .Y(_218_) );
NOR2X1 NOR2X1_84 ( .A(reset_bF_buf4), .B(_218_), .Y(keyreg1__3__3_) );
DFFPOSX1 DFFPOSX1_119 ( .CLK(reset_bF_buf3), .D(keyreg1__0__0_), .Q(alreg1_new_alarm_ls_hr_0_) );
DFFPOSX1 DFFPOSX1_120 ( .CLK(reset_bF_buf2), .D(keyreg1__0__1_), .Q(alreg1_new_alarm_ls_hr_1_) );
DFFPOSX1 DFFPOSX1_121 ( .CLK(reset_bF_buf1), .D(keyreg1__0__2_), .Q(alreg1_new_alarm_ls_hr_2_) );
DFFPOSX1 DFFPOSX1_122 ( .CLK(reset_bF_buf0), .D(keyreg1__0__3_), .Q(alreg1_new_alarm_ls_hr_3_) );
DFFPOSX1 DFFPOSX1_123 ( .CLK(reset_bF_buf9), .D(keyreg1__1__0_), .Q(alreg1_new_alarm_ls_min_0_) );
DFFPOSX1 DFFPOSX1_124 ( .CLK(reset_bF_buf8), .D(keyreg1__1__1_), .Q(alreg1_new_alarm_ls_min_1_) );
DFFPOSX1 DFFPOSX1_125 ( .CLK(reset_bF_buf7), .D(keyreg1__1__2_), .Q(alreg1_new_alarm_ls_min_2_) );
DFFPOSX1 DFFPOSX1_126 ( .CLK(reset_bF_buf6), .D(keyreg1__1__3_), .Q(alreg1_new_alarm_ls_min_3_) );
DFFPOSX1 DFFPOSX1_127 ( .CLK(reset_bF_buf5), .D(keyreg1__2__0_), .Q(alreg1_new_alarm_ms_hr_0_) );
DFFPOSX1 DFFPOSX1_128 ( .CLK(reset_bF_buf4), .D(keyreg1__2__1_), .Q(alreg1_new_alarm_ms_hr_1_) );
DFFPOSX1 DFFPOSX1_129 ( .CLK(reset_bF_buf3), .D(keyreg1__2__2_), .Q(alreg1_new_alarm_ms_hr_2_) );
DFFPOSX1 DFFPOSX1_130 ( .CLK(reset_bF_buf2), .D(keyreg1__2__3_), .Q(alreg1_new_alarm_ms_hr_3_) );
DFFPOSX1 DFFPOSX1_131 ( .CLK(reset_bF_buf1), .D(keyreg1__3__0_), .Q(alreg1_new_alarm_ms_min_0_) );
DFFPOSX1 DFFPOSX1_132 ( .CLK(reset_bF_buf0), .D(keyreg1__3__1_), .Q(alreg1_new_alarm_ms_min_1_) );
DFFPOSX1 DFFPOSX1_133 ( .CLK(reset_bF_buf9), .D(keyreg1__3__2_), .Q(alreg1_new_alarm_ms_min_2_) );
DFFPOSX1 DFFPOSX1_134 ( .CLK(reset_bF_buf8), .D(keyreg1__3__3_), .Q(alreg1_new_alarm_ms_min_3_) );
DFFPOSX1 DFFPOSX1_135 ( .CLK(clock_bF_buf4), .D(keyreg1__0__0_), .Q(alreg1_new_alarm_ls_hr_0_) );
DFFPOSX1 DFFPOSX1_136 ( .CLK(clock_bF_buf3), .D(keyreg1__0__1_), .Q(alreg1_new_alarm_ls_hr_1_) );
DFFPOSX1 DFFPOSX1_137 ( .CLK(clock_bF_buf2), .D(keyreg1__0__2_), .Q(alreg1_new_alarm_ls_hr_2_) );
DFFPOSX1 DFFPOSX1_138 ( .CLK(clock_bF_buf1), .D(keyreg1__0__3_), .Q(alreg1_new_alarm_ls_hr_3_) );
DFFPOSX1 DFFPOSX1_139 ( .CLK(clock_bF_buf0), .D(keyreg1__1__0_), .Q(alreg1_new_alarm_ls_min_0_) );
DFFPOSX1 DFFPOSX1_140 ( .CLK(clock_bF_buf7), .D(keyreg1__1__1_), .Q(alreg1_new_alarm_ls_min_1_) );
DFFPOSX1 DFFPOSX1_141 ( .CLK(clock_bF_buf6), .D(keyreg1__1__2_), .Q(alreg1_new_alarm_ls_min_2_) );
DFFPOSX1 DFFPOSX1_142 ( .CLK(clock_bF_buf5), .D(keyreg1__1__3_), .Q(alreg1_new_alarm_ls_min_3_) );
DFFPOSX1 DFFPOSX1_143 ( .CLK(clock_bF_buf4), .D(keyreg1__2__0_), .Q(alreg1_new_alarm_ms_hr_0_) );
DFFPOSX1 DFFPOSX1_144 ( .CLK(clock_bF_buf3), .D(keyreg1__2__1_), .Q(alreg1_new_alarm_ms_hr_1_) );
DFFPOSX1 DFFPOSX1_145 ( .CLK(clock_bF_buf2), .D(keyreg1__2__2_), .Q(alreg1_new_alarm_ms_hr_2_) );
DFFPOSX1 DFFPOSX1_146 ( .CLK(clock_bF_buf1), .D(keyreg1__2__3_), .Q(alreg1_new_alarm_ms_hr_3_) );
DFFPOSX1 DFFPOSX1_147 ( .CLK(clock_bF_buf0), .D(keyreg1__3__0_), .Q(alreg1_new_alarm_ms_min_0_) );
DFFPOSX1 DFFPOSX1_148 ( .CLK(clock_bF_buf7), .D(keyreg1__3__1_), .Q(alreg1_new_alarm_ms_min_1_) );
DFFPOSX1 DFFPOSX1_149 ( .CLK(clock_bF_buf6), .D(keyreg1__3__2_), .Q(alreg1_new_alarm_ms_min_2_) );
DFFPOSX1 DFFPOSX1_150 ( .CLK(clock_bF_buf5), .D(keyreg1__3__3_), .Q(alreg1_new_alarm_ms_min_3_) );
NAND2X1 NAND2X1_32 ( .A(lcd_disp_LS_HR_sound_alarm), .B(lcd_disp_MS_HR_sound_alarm), .Y(_219_) );
NAND2X1 NAND2X1_33 ( .A(lcd_disp_MS_MIN_sound_alarm), .B(lcd_disp_LS_MIN_sound_alarm), .Y(_220_) );
NOR2X1 NOR2X1_85 ( .A(_219_), .B(_220_), .Y(_0_) );
NOR2X1 NOR2X1_86 ( .A(alarm_time_ls_hr_0_), .B(count1_current_time_ls_hr_0_), .Y(_223_) );
AND2X2 AND2X2_11 ( .A(alarm_time_ls_hr_0_), .B(count1_current_time_ls_hr_0_), .Y(_224_) );
AND2X2 AND2X2_12 ( .A(alarm_time_ls_hr_1_), .B(count1_current_time_ls_hr_1_), .Y(_225_) );
NOR2X1 NOR2X1_87 ( .A(alarm_time_ls_hr_1_), .B(count1_current_time_ls_hr_1_), .Y(_226_) );
OAI22X1 OAI22X1_1 ( .A(_224_), .B(_223_), .C(_225_), .D(_226_), .Y(_227_) );
XOR2X1 XOR2X1_1 ( .A(alarm_time_ls_hr_3_), .B(count1_current_time_ls_hr_3_), .Y(_228_) );
XOR2X1 XOR2X1_2 ( .A(alarm_time_ls_hr_2_), .B(count1_current_time_ls_hr_2_), .Y(_229_) );
NOR3X1 NOR3X1_9 ( .A(_228_), .B(_229_), .C(_227_), .Y(lcd_disp_LS_HR_sound_alarm) );
INVX1 INVX1_35 ( .A(count1_current_time_ls_hr_0_), .Y(_230_) );
NAND2X1 NAND2X1_34 ( .A(alarm_time_ls_hr_0_), .B(fsm1__25__bF_buf3), .Y(_231_) );
OAI21X1 OAI21X1_46 ( .A(_230_), .B(fsm1__25__bF_buf2), .C(_231_), .Y(_221__0_) );
INVX1 INVX1_36 ( .A(count1_current_time_ls_hr_1_), .Y(_232_) );
NAND2X1 NAND2X1_35 ( .A(alarm_time_ls_hr_1_), .B(fsm1__25__bF_buf1), .Y(_233_) );
OAI21X1 OAI21X1_47 ( .A(_232_), .B(fsm1__25__bF_buf0), .C(_233_), .Y(_221__1_) );
INVX1 INVX1_37 ( .A(count1_current_time_ls_hr_2_), .Y(_234_) );
NAND2X1 NAND2X1_36 ( .A(alarm_time_ls_hr_2_), .B(fsm1__25__bF_buf4), .Y(_235_) );
OAI21X1 OAI21X1_48 ( .A(_234_), .B(fsm1__25__bF_buf3), .C(_235_), .Y(_221__2_) );
INVX1 INVX1_38 ( .A(count1_current_time_ls_hr_3_), .Y(_236_) );
NAND2X1 NAND2X1_37 ( .A(alarm_time_ls_hr_3_), .B(fsm1__25__bF_buf2), .Y(_237_) );
OAI21X1 OAI21X1_49 ( .A(_236_), .B(fsm1__25__bF_buf1), .C(_237_), .Y(_221__3_) );
MUX2X1 MUX2X1_33 ( .A(alreg1_new_alarm_ls_hr_0_), .B(lcd_disp_LS_HR__6__0_), .S(fsm1_show_new_time_bF_buf3), .Y(_238_) );
MUX2X1 MUX2X1_34 ( .A(alreg1_new_alarm_ls_hr_3_), .B(lcd_disp_LS_HR__6__3_), .S(fsm1_show_new_time_bF_buf2), .Y(_239_) );
MUX2X1 MUX2X1_35 ( .A(alreg1_new_alarm_ls_hr_1_), .B(lcd_disp_LS_HR__6__1_), .S(fsm1_show_new_time_bF_buf1), .Y(_240_) );
MUX2X1 MUX2X1_36 ( .A(alreg1_new_alarm_ls_hr_2_), .B(lcd_disp_LS_HR__6__2_), .S(fsm1_show_new_time_bF_buf0), .Y(_241_) );
AOI21X1 AOI21X1_33 ( .A(_240_), .B(_241_), .C(_239_), .Y(_242_) );
NOR2X1 NOR2X1_88 ( .A(_238_), .B(_242_), .Y(_1__0_) );
OAI21X1 OAI21X1_50 ( .A(_239_), .B(_241_), .C(_240_), .Y(_1__1_) );
INVX1 INVX1_39 ( .A(_239_), .Y(_1__3_) );
NOR2X1 NOR2X1_89 ( .A(_241_), .B(_1__3_), .Y(_1__2_) );
INVX1 INVX1_40 ( .A(fsm1_show_new_time_bF_buf3), .Y(_222_) );
NOR2X1 NOR2X1_90 ( .A(alarm_time_ls_min_0_), .B(count1_current_time_ls_min_0_), .Y(_245_) );
AND2X2 AND2X2_13 ( .A(alarm_time_ls_min_0_), .B(count1_current_time_ls_min_0_), .Y(_246_) );
AND2X2 AND2X2_14 ( .A(alarm_time_ls_min_1_), .B(count1_current_time_ls_min_1_), .Y(_247_) );
NOR2X1 NOR2X1_91 ( .A(alarm_time_ls_min_1_), .B(count1_current_time_ls_min_1_), .Y(_248_) );
OAI22X1 OAI22X1_2 ( .A(_246_), .B(_245_), .C(_247_), .D(_248_), .Y(_249_) );
XOR2X1 XOR2X1_3 ( .A(alarm_time_ls_min_3_), .B(count1_current_time_ls_min_3_), .Y(_250_) );
XOR2X1 XOR2X1_4 ( .A(alarm_time_ls_min_2_), .B(count1_current_time_ls_min_2_), .Y(_251_) );
NOR3X1 NOR3X1_10 ( .A(_250_), .B(_251_), .C(_249_), .Y(lcd_disp_LS_MIN_sound_alarm) );
INVX1 INVX1_41 ( .A(count1_current_time_ls_min_0_), .Y(_252_) );
NAND2X1 NAND2X1_38 ( .A(alarm_time_ls_min_0_), .B(fsm1__25__bF_buf0), .Y(_253_) );
OAI21X1 OAI21X1_51 ( .A(_252_), .B(fsm1__25__bF_buf4), .C(_253_), .Y(_243__0_) );
INVX1 INVX1_42 ( .A(count1_current_time_ls_min_1_), .Y(_254_) );
NAND2X1 NAND2X1_39 ( .A(alarm_time_ls_min_1_), .B(fsm1__25__bF_buf3), .Y(_255_) );
OAI21X1 OAI21X1_52 ( .A(_254_), .B(fsm1__25__bF_buf2), .C(_255_), .Y(_243__1_) );
INVX1 INVX1_43 ( .A(count1_current_time_ls_min_2_), .Y(_256_) );
NAND2X1 NAND2X1_40 ( .A(alarm_time_ls_min_2_), .B(fsm1__25__bF_buf1), .Y(_257_) );
OAI21X1 OAI21X1_53 ( .A(_256_), .B(fsm1__25__bF_buf0), .C(_257_), .Y(_243__2_) );
INVX1 INVX1_44 ( .A(count1_current_time_ls_min_3_), .Y(_258_) );
NAND2X1 NAND2X1_41 ( .A(alarm_time_ls_min_3_), .B(fsm1__25__bF_buf4), .Y(_259_) );
OAI21X1 OAI21X1_54 ( .A(_258_), .B(fsm1__25__bF_buf3), .C(_259_), .Y(_243__3_) );
MUX2X1 MUX2X1_37 ( .A(alreg1_new_alarm_ls_min_0_), .B(lcd_disp_LS_MIN__6__0_), .S(fsm1_show_new_time_bF_buf2), .Y(_260_) );
MUX2X1 MUX2X1_38 ( .A(alreg1_new_alarm_ls_min_3_), .B(lcd_disp_LS_MIN__6__3_), .S(fsm1_show_new_time_bF_buf1), .Y(_261_) );
MUX2X1 MUX2X1_39 ( .A(alreg1_new_alarm_ls_min_1_), .B(lcd_disp_LS_MIN__6__1_), .S(fsm1_show_new_time_bF_buf0), .Y(_262_) );
MUX2X1 MUX2X1_40 ( .A(alreg1_new_alarm_ls_min_2_), .B(lcd_disp_LS_MIN__6__2_), .S(fsm1_show_new_time_bF_buf3), .Y(_263_) );
AOI21X1 AOI21X1_34 ( .A(_262_), .B(_263_), .C(_261_), .Y(_264_) );
NOR2X1 NOR2X1_92 ( .A(_260_), .B(_264_), .Y(_2__0_) );
OAI21X1 OAI21X1_55 ( .A(_261_), .B(_263_), .C(_262_), .Y(_2__1_) );
INVX1 INVX1_45 ( .A(_261_), .Y(_2__3_) );
NOR2X1 NOR2X1_93 ( .A(_263_), .B(_2__3_), .Y(_2__2_) );
INVX1 INVX1_46 ( .A(fsm1_show_new_time_bF_buf2), .Y(_244_) );
NOR2X1 NOR2X1_94 ( .A(alarm_time_ms_hr_0_), .B(count1_current_time_ms_hr_0_), .Y(_267_) );
AND2X2 AND2X2_15 ( .A(alarm_time_ms_hr_0_), .B(count1_current_time_ms_hr_0_), .Y(_268_) );
AND2X2 AND2X2_16 ( .A(alarm_time_ms_hr_1_), .B(count1_current_time_ms_hr_1_), .Y(_269_) );
NOR2X1 NOR2X1_95 ( .A(alarm_time_ms_hr_1_), .B(count1_current_time_ms_hr_1_), .Y(_270_) );
OAI22X1 OAI22X1_3 ( .A(_268_), .B(_267_), .C(_269_), .D(_270_), .Y(_271_) );
XOR2X1 XOR2X1_5 ( .A(alarm_time_ms_hr_3_), .B(count1_current_time_ms_hr_3_), .Y(_272_) );
XOR2X1 XOR2X1_6 ( .A(alarm_time_ms_hr_2_), .B(count1_current_time_ms_hr_2_), .Y(_273_) );
NOR3X1 NOR3X1_11 ( .A(_272_), .B(_273_), .C(_271_), .Y(lcd_disp_MS_HR_sound_alarm) );
INVX1 INVX1_47 ( .A(count1_current_time_ms_hr_0_), .Y(_274_) );
NAND2X1 NAND2X1_42 ( .A(alarm_time_ms_hr_0_), .B(fsm1__25__bF_buf2), .Y(_275_) );
OAI21X1 OAI21X1_56 ( .A(_274_), .B(fsm1__25__bF_buf1), .C(_275_), .Y(_265__0_) );
INVX1 INVX1_48 ( .A(count1_current_time_ms_hr_1_), .Y(_276_) );
NAND2X1 NAND2X1_43 ( .A(alarm_time_ms_hr_1_), .B(fsm1__25__bF_buf0), .Y(_277_) );
OAI21X1 OAI21X1_57 ( .A(_276_), .B(fsm1__25__bF_buf4), .C(_277_), .Y(_265__1_) );
INVX1 INVX1_49 ( .A(count1_current_time_ms_hr_2_), .Y(_278_) );
NAND2X1 NAND2X1_44 ( .A(alarm_time_ms_hr_2_), .B(fsm1__25__bF_buf3), .Y(_279_) );
OAI21X1 OAI21X1_58 ( .A(_278_), .B(fsm1__25__bF_buf2), .C(_279_), .Y(_265__2_) );
INVX1 INVX1_50 ( .A(count1_current_time_ms_hr_3_), .Y(_280_) );
NAND2X1 NAND2X1_45 ( .A(alarm_time_ms_hr_3_), .B(fsm1__25__bF_buf1), .Y(_281_) );
OAI21X1 OAI21X1_59 ( .A(_280_), .B(fsm1__25__bF_buf0), .C(_281_), .Y(_265__3_) );
MUX2X1 MUX2X1_41 ( .A(alreg1_new_alarm_ms_hr_0_), .B(lcd_disp_MS_HR__6__0_), .S(fsm1_show_new_time_bF_buf1), .Y(_282_) );
MUX2X1 MUX2X1_42 ( .A(alreg1_new_alarm_ms_hr_3_), .B(lcd_disp_MS_HR__6__3_), .S(fsm1_show_new_time_bF_buf0), .Y(_283_) );
MUX2X1 MUX2X1_43 ( .A(alreg1_new_alarm_ms_hr_1_), .B(lcd_disp_MS_HR__6__1_), .S(fsm1_show_new_time_bF_buf3), .Y(_284_) );
MUX2X1 MUX2X1_44 ( .A(alreg1_new_alarm_ms_hr_2_), .B(lcd_disp_MS_HR__6__2_), .S(fsm1_show_new_time_bF_buf2), .Y(_285_) );
AOI21X1 AOI21X1_35 ( .A(_284_), .B(_285_), .C(_283_), .Y(_286_) );
NOR2X1 NOR2X1_96 ( .A(_282_), .B(_286_), .Y(_3__0_) );
OAI21X1 OAI21X1_60 ( .A(_283_), .B(_285_), .C(_284_), .Y(_3__1_) );
INVX1 INVX1_51 ( .A(_283_), .Y(_3__3_) );
NOR2X1 NOR2X1_97 ( .A(_285_), .B(_3__3_), .Y(_3__2_) );
INVX1 INVX1_52 ( .A(fsm1_show_new_time_bF_buf1), .Y(_266_) );
NOR2X1 NOR2X1_98 ( .A(alarm_time_ms_min_0_), .B(count1_current_time_ms_min_0_), .Y(_289_) );
AND2X2 AND2X2_17 ( .A(alarm_time_ms_min_0_), .B(count1_current_time_ms_min_0_), .Y(_290_) );
AND2X2 AND2X2_18 ( .A(alarm_time_ms_min_1_), .B(count1_current_time_ms_min_1_), .Y(_291_) );
NOR2X1 NOR2X1_99 ( .A(alarm_time_ms_min_1_), .B(count1_current_time_ms_min_1_), .Y(_292_) );
OAI22X1 OAI22X1_4 ( .A(_290_), .B(_289_), .C(_291_), .D(_292_), .Y(_293_) );
XOR2X1 XOR2X1_7 ( .A(alarm_time_ms_min_3_), .B(count1_current_time_ms_min_3_), .Y(_294_) );
XOR2X1 XOR2X1_8 ( .A(alarm_time_ms_min_2_), .B(count1_current_time_ms_min_2_), .Y(_295_) );
NOR3X1 NOR3X1_12 ( .A(_294_), .B(_295_), .C(_293_), .Y(lcd_disp_MS_MIN_sound_alarm) );
INVX1 INVX1_53 ( .A(count1_current_time_ms_min_0_), .Y(_296_) );
NAND2X1 NAND2X1_46 ( .A(alarm_time_ms_min_0_), .B(fsm1__25__bF_buf4), .Y(_297_) );
OAI21X1 OAI21X1_61 ( .A(_296_), .B(fsm1__25__bF_buf3), .C(_297_), .Y(_287__0_) );
INVX1 INVX1_54 ( .A(count1_current_time_ms_min_1_), .Y(_298_) );
NAND2X1 NAND2X1_47 ( .A(alarm_time_ms_min_1_), .B(fsm1__25__bF_buf2), .Y(_299_) );
OAI21X1 OAI21X1_62 ( .A(_298_), .B(fsm1__25__bF_buf1), .C(_299_), .Y(_287__1_) );
INVX1 INVX1_55 ( .A(count1_current_time_ms_min_2_), .Y(_300_) );
NAND2X1 NAND2X1_48 ( .A(alarm_time_ms_min_2_), .B(fsm1__25__bF_buf0), .Y(_301_) );
OAI21X1 OAI21X1_63 ( .A(_300_), .B(fsm1__25__bF_buf4), .C(_301_), .Y(_287__2_) );
INVX1 INVX1_56 ( .A(count1_current_time_ms_min_3_), .Y(_302_) );
NAND2X1 NAND2X1_49 ( .A(alarm_time_ms_min_3_), .B(fsm1__25__bF_buf3), .Y(_303_) );
OAI21X1 OAI21X1_64 ( .A(_302_), .B(fsm1__25__bF_buf2), .C(_303_), .Y(_287__3_) );
MUX2X1 MUX2X1_45 ( .A(alreg1_new_alarm_ms_min_0_), .B(lcd_disp_MS_MIN__6__0_), .S(fsm1_show_new_time_bF_buf0), .Y(_304_) );
MUX2X1 MUX2X1_46 ( .A(alreg1_new_alarm_ms_min_3_), .B(lcd_disp_MS_MIN__6__3_), .S(fsm1_show_new_time_bF_buf3), .Y(_305_) );
MUX2X1 MUX2X1_47 ( .A(alreg1_new_alarm_ms_min_1_), .B(lcd_disp_MS_MIN__6__1_), .S(fsm1_show_new_time_bF_buf2), .Y(_306_) );
MUX2X1 MUX2X1_48 ( .A(alreg1_new_alarm_ms_min_2_), .B(lcd_disp_MS_MIN__6__2_), .S(fsm1_show_new_time_bF_buf1), .Y(_307_) );
AOI21X1 AOI21X1_36 ( .A(_306_), .B(_307_), .C(_305_), .Y(_308_) );
NOR2X1 NOR2X1_100 ( .A(_304_), .B(_308_), .Y(_4__0_) );
OAI21X1 OAI21X1_65 ( .A(_305_), .B(_307_), .C(_306_), .Y(_4__1_) );
INVX1 INVX1_57 ( .A(_305_), .Y(_4__3_) );
NOR2X1 NOR2X1_101 ( .A(_307_), .B(_4__3_), .Y(_4__2_) );
INVX1 INVX1_58 ( .A(fsm1_show_new_time_bF_buf0), .Y(_288_) );
NAND2X1 NAND2X1_50 ( .A(tgen1_count_4_), .B(tgen1_count_7_), .Y(_317_) );
NAND2X1 NAND2X1_51 ( .A(tgen1_count_5_), .B(tgen1_count_6_), .Y(_318_) );
NOR2X1 NOR2X1_102 ( .A(_317_), .B(_318_), .Y(_319_) );
NAND2X1 NAND2X1_52 ( .A(tgen1_count_0_), .B(tgen1_count_1_), .Y(_320_) );
NAND2X1 NAND2X1_53 ( .A(tgen1_count_3_), .B(tgen1_count_2_), .Y(_321_) );
NOR2X1 NOR2X1_103 ( .A(_320_), .B(_321_), .Y(_322_) );
NAND2X1 NAND2X1_54 ( .A(_319_), .B(_322_), .Y(_323_) );
NOR2X1 NOR2X1_104 ( .A(reset_bF_buf7), .B(count1_load_new_c), .Y(_324_) );
INVX2 INVX2_15 ( .A(_324_), .Y(_325_) );
NOR2X1 NOR2X1_105 ( .A(_325_), .B(_323_), .Y(tgen1__03_) );
INVX1 INVX1_59 ( .A(tgen1_one_minute_reg), .Y(_326_) );
NAND2X1 NAND2X1_55 ( .A(fsm1_one_second), .B(fastwatch), .Y(_327_) );
OAI21X1 OAI21X1_66 ( .A(_326_), .B(fastwatch), .C(_327_), .Y(count1_one_minute) );
AND2X2 AND2X2_19 ( .A(tgen1_count_4_), .B(tgen1_count_7_), .Y(_328_) );
AND2X2 AND2X2_20 ( .A(tgen1_count_5_), .B(tgen1_count_6_), .Y(_329_) );
NAND2X1 NAND2X1_56 ( .A(_328_), .B(_329_), .Y(_330_) );
OR2X2 OR2X2_10 ( .A(_320_), .B(_321_), .Y(_331_) );
NAND2X1 NAND2X1_57 ( .A(tgen1_count_9_), .B(tgen1_count_8_), .Y(_332_) );
NOR3X1 NOR3X1_13 ( .A(_330_), .B(_332_), .C(_331_), .Y(_333_) );
NAND2X1 NAND2X1_58 ( .A(tgen1_count_11_), .B(tgen1_count_12_), .Y(_334_) );
INVX2 INVX2_16 ( .A(tgen1_count_10_), .Y(_335_) );
NAND2X1 NAND2X1_59 ( .A(tgen1_count_13_), .B(_335_), .Y(_336_) );
NOR2X1 NOR2X1_106 ( .A(_334_), .B(_336_), .Y(_337_) );
NAND2X1 NAND2X1_60 ( .A(_337_), .B(_333_), .Y(_338_) );
NOR2X1 NOR2X1_107 ( .A(_325_), .B(_338_), .Y(tgen1__02_) );
NOR2X1 NOR2X1_108 ( .A(tgen1_count_0_), .B(_325_), .Y(tgen1__00__0_) );
INVX2 INVX2_17 ( .A(_320_), .Y(_339_) );
OAI21X1 OAI21X1_67 ( .A(tgen1_count_0_), .B(tgen1_count_1_), .C(_324_), .Y(_340_) );
NOR2X1 NOR2X1_109 ( .A(_339_), .B(_340_), .Y(tgen1__00__1_) );
OAI21X1 OAI21X1_68 ( .A(_339_), .B(tgen1_count_2_), .C(_324_), .Y(_341_) );
BUFX2 BUFX2_34 ( .A(1'b1), .Y(_1__4_) );
BUFX2 BUFX2_35 ( .A(1'b1), .Y(_1__5_) );
BUFX2 BUFX2_36 ( .A(1'b0), .Y(_1__6_) );
BUFX2 BUFX2_37 ( .A(1'b0), .Y(_1__7_) );
BUFX2 BUFX2_38 ( .A(1'b1), .Y(_2__4_) );
BUFX2 BUFX2_39 ( .A(1'b1), .Y(_2__5_) );
BUFX2 BUFX2_40 ( .A(1'b0), .Y(_2__6_) );
BUFX2 BUFX2_41 ( .A(1'b0), .Y(_2__7_) );
BUFX2 BUFX2_42 ( .A(1'b1), .Y(_3__4_) );
BUFX2 BUFX2_43 ( .A(1'b1), .Y(_3__5_) );
BUFX2 BUFX2_44 ( .A(1'b0), .Y(_3__6_) );
BUFX2 BUFX2_45 ( .A(1'b0), .Y(_3__7_) );
BUFX2 BUFX2_46 ( .A(1'b1), .Y(_4__4_) );
BUFX2 BUFX2_47 ( .A(1'b1), .Y(_4__5_) );
BUFX2 BUFX2_48 ( .A(1'b0), .Y(_4__6_) );
BUFX2 BUFX2_49 ( .A(1'b0), .Y(_4__7_) );
BUFX2 BUFX2_50 ( .A(_127__2_), .Y(_127__1_) );
BUFX2 BUFX2_51 ( .A(1'b0), .Y(_128__0_) );
BUFX2 BUFX2_52 ( .A(_128__2_), .Y(_128__1_) );
BUFX2 BUFX2_53 ( .A(fsm1__04__1_), .Y(fsm1__04__0_) );
BUFX2 BUFX2_54 ( .A(fsm1__07__2_), .Y(fsm1__07__0_) );
BUFX2 BUFX2_55 ( .A(fsm1__08__2_), .Y(fsm1__08__1_) );
BUFX2 BUFX2_56 ( .A(fsm1__09__2_), .Y(fsm1__09__1_) );
endmodule
