VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO alarm_clock_top
  CLASS BLOCK ;
  FOREIGN alarm_clock_top ;
  ORIGIN 2.600 3.000 ;
  SIZE 201.200 BY 176.200 ;
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT 132.600 166.100 133.000 166.600 ;
        RECT 133.400 166.100 133.800 166.600 ;
        RECT 132.600 165.800 133.800 166.100 ;
        RECT 173.400 165.800 173.800 166.600 ;
        RECT 187.800 165.800 188.200 166.600 ;
        RECT 190.200 165.800 190.600 166.600 ;
        RECT 1.400 160.800 1.800 164.500 ;
        RECT 3.800 160.800 4.200 164.500 ;
        RECT 7.000 160.800 7.400 165.100 ;
        RECT 8.600 160.800 9.000 163.100 ;
        RECT 9.400 160.800 9.800 165.100 ;
        RECT 11.500 160.800 11.900 163.100 ;
        RECT 14.200 160.800 14.600 164.500 ;
        RECT 16.600 160.800 17.000 164.500 ;
        RECT 19.800 160.800 20.200 165.100 ;
        RECT 21.400 160.800 21.800 164.500 ;
        RECT 23.800 160.800 24.200 165.100 ;
        RECT 26.600 160.800 27.000 163.100 ;
        RECT 28.200 160.800 28.600 163.100 ;
        RECT 31.000 160.800 31.400 165.000 ;
        RECT 33.400 160.800 33.800 165.100 ;
        RECT 36.200 160.800 36.600 163.100 ;
        RECT 37.800 160.800 38.200 163.100 ;
        RECT 40.600 160.800 41.000 165.000 ;
        RECT 42.200 160.800 42.600 165.100 ;
        RECT 47.000 160.800 47.400 164.900 ;
        RECT 49.600 160.800 50.000 165.100 ;
        RECT 51.800 160.800 52.200 165.100 ;
        RECT 54.600 160.800 55.000 163.100 ;
        RECT 56.200 160.800 56.600 163.100 ;
        RECT 59.000 160.800 59.400 165.000 ;
        RECT 62.200 160.800 62.600 165.100 ;
        RECT 63.800 160.800 64.200 165.100 ;
        RECT 66.600 160.800 67.000 163.100 ;
        RECT 68.200 160.800 68.600 163.100 ;
        RECT 71.000 160.800 71.400 165.000 ;
        RECT 73.400 160.800 73.800 165.100 ;
        RECT 76.200 160.800 76.600 163.100 ;
        RECT 77.800 160.800 78.200 163.100 ;
        RECT 80.600 160.800 81.000 165.000 ;
        RECT 83.000 160.800 83.400 164.500 ;
        RECT 84.600 160.800 85.000 165.100 ;
        RECT 87.800 160.800 88.200 164.500 ;
        RECT 90.200 160.800 90.600 163.100 ;
        RECT 91.800 160.800 92.200 165.100 ;
        RECT 94.600 160.800 95.000 163.100 ;
        RECT 96.200 160.800 96.600 163.100 ;
        RECT 99.000 160.800 99.400 165.000 ;
        RECT 102.200 160.800 102.600 165.100 ;
        RECT 105.400 160.800 105.800 164.500 ;
        RECT 107.800 160.800 108.200 165.100 ;
        RECT 110.600 160.800 111.000 163.100 ;
        RECT 112.200 160.800 112.600 163.100 ;
        RECT 115.000 160.800 115.400 165.000 ;
        RECT 117.400 160.800 117.800 164.500 ;
        RECT 119.800 160.800 120.200 164.500 ;
        RECT 122.200 160.800 122.600 165.100 ;
        RECT 125.000 160.800 125.400 163.100 ;
        RECT 126.600 160.800 127.000 163.100 ;
        RECT 129.400 160.800 129.800 165.000 ;
        RECT 131.800 160.800 132.200 164.500 ;
        RECT 134.200 160.800 134.600 164.500 ;
        RECT 136.600 160.800 137.000 165.000 ;
        RECT 139.400 160.800 139.800 163.100 ;
        RECT 141.000 160.800 141.400 163.100 ;
        RECT 143.800 160.800 144.200 165.100 ;
        RECT 145.400 160.800 145.800 165.100 ;
        RECT 150.200 160.800 150.600 164.900 ;
        RECT 152.800 160.800 153.200 165.100 ;
        RECT 155.000 160.800 155.400 165.100 ;
        RECT 157.800 160.800 158.200 163.100 ;
        RECT 159.400 160.800 159.800 163.100 ;
        RECT 162.200 160.800 162.600 165.000 ;
        RECT 164.600 160.800 165.000 165.000 ;
        RECT 167.400 160.800 167.800 163.100 ;
        RECT 169.000 160.800 169.400 163.100 ;
        RECT 171.800 160.800 172.200 165.100 ;
        RECT 174.200 160.800 174.600 164.500 ;
        RECT 176.600 160.800 177.000 165.100 ;
        RECT 179.400 160.800 179.800 163.100 ;
        RECT 181.000 160.800 181.400 163.100 ;
        RECT 183.800 160.800 184.200 165.000 ;
        RECT 186.200 160.800 186.600 164.500 ;
        RECT 188.600 160.800 189.000 164.500 ;
        RECT 191.000 160.800 191.400 164.500 ;
        RECT 192.600 160.800 193.000 163.100 ;
        RECT 0.200 160.200 195.800 160.800 ;
        RECT 1.400 155.900 1.800 160.200 ;
        RECT 4.200 157.900 4.600 160.200 ;
        RECT 5.800 157.900 6.200 160.200 ;
        RECT 8.600 156.000 9.000 160.200 ;
        RECT 10.800 155.900 11.200 160.200 ;
        RECT 13.400 156.100 13.800 160.200 ;
        RECT 15.600 155.900 16.000 160.200 ;
        RECT 18.200 156.100 18.600 160.200 ;
        RECT 20.400 155.900 20.800 160.200 ;
        RECT 23.000 156.100 23.400 160.200 ;
        RECT 25.200 155.900 25.600 160.200 ;
        RECT 27.800 156.100 28.200 160.200 ;
        RECT 30.200 155.900 30.600 160.200 ;
        RECT 33.000 157.900 33.400 160.200 ;
        RECT 34.600 157.900 35.000 160.200 ;
        RECT 37.400 156.000 37.800 160.200 ;
        RECT 39.800 156.000 40.200 160.200 ;
        RECT 42.600 157.900 43.000 160.200 ;
        RECT 44.200 157.900 44.600 160.200 ;
        RECT 47.000 155.900 47.400 160.200 ;
        RECT 51.000 157.900 51.400 160.200 ;
        RECT 52.600 155.900 53.000 160.200 ;
        RECT 55.400 157.900 55.800 160.200 ;
        RECT 57.000 157.900 57.400 160.200 ;
        RECT 59.800 156.000 60.200 160.200 ;
        RECT 62.200 155.900 62.600 160.200 ;
        RECT 65.000 157.900 65.400 160.200 ;
        RECT 66.600 157.900 67.000 160.200 ;
        RECT 69.400 156.000 69.800 160.200 ;
        RECT 71.800 155.900 72.200 160.200 ;
        RECT 74.600 157.900 75.000 160.200 ;
        RECT 76.200 157.900 76.600 160.200 ;
        RECT 79.000 156.000 79.400 160.200 ;
        RECT 81.400 155.900 81.800 160.200 ;
        RECT 84.200 157.900 84.600 160.200 ;
        RECT 85.800 157.900 86.200 160.200 ;
        RECT 88.600 156.000 89.000 160.200 ;
        RECT 90.800 155.900 91.200 160.200 ;
        RECT 93.400 156.100 93.800 160.200 ;
        RECT 95.800 156.500 96.200 160.200 ;
        RECT 99.800 155.900 100.200 160.200 ;
        RECT 101.900 157.900 102.300 160.200 ;
        RECT 104.600 155.900 105.000 160.200 ;
        RECT 106.200 156.500 106.600 160.200 ;
        RECT 108.600 156.500 109.000 160.200 ;
        RECT 111.000 156.100 111.400 160.200 ;
        RECT 113.600 155.900 114.000 160.200 ;
        RECT 115.800 156.500 116.200 160.200 ;
        RECT 117.400 155.900 117.800 160.200 ;
        RECT 121.400 156.500 121.800 160.200 ;
        RECT 123.300 157.900 123.700 160.200 ;
        RECT 125.400 155.900 125.800 160.200 ;
        RECT 126.200 157.900 126.600 160.200 ;
        RECT 127.800 155.900 128.200 160.200 ;
        RECT 131.000 156.500 131.400 160.200 ;
        RECT 134.200 155.900 134.600 160.200 ;
        RECT 135.800 155.900 136.200 160.200 ;
        RECT 138.600 157.900 139.000 160.200 ;
        RECT 140.200 157.900 140.600 160.200 ;
        RECT 143.000 156.000 143.400 160.200 ;
        RECT 145.200 155.900 145.600 160.200 ;
        RECT 147.800 156.100 148.200 160.200 ;
        RECT 152.600 155.900 153.000 160.200 ;
        RECT 154.200 156.000 154.600 160.200 ;
        RECT 157.000 157.900 157.400 160.200 ;
        RECT 158.600 157.900 159.000 160.200 ;
        RECT 161.400 155.900 161.800 160.200 ;
        RECT 163.800 156.100 164.200 160.200 ;
        RECT 165.400 157.900 165.800 160.200 ;
        RECT 166.200 155.900 166.600 160.200 ;
        RECT 169.200 155.900 169.600 160.200 ;
        RECT 171.800 156.100 172.200 160.200 ;
        RECT 174.200 156.100 174.600 160.200 ;
        RECT 176.800 155.900 177.200 160.200 ;
        RECT 179.000 156.500 179.400 160.200 ;
        RECT 182.200 155.900 182.600 160.200 ;
        RECT 183.800 156.000 184.200 160.200 ;
        RECT 186.600 157.900 187.000 160.200 ;
        RECT 188.200 157.900 188.600 160.200 ;
        RECT 191.000 155.900 191.400 160.200 ;
        RECT 193.400 156.500 193.800 160.200 ;
        RECT 179.800 154.400 180.200 155.200 ;
        RECT 192.600 154.400 193.000 155.200 ;
        RECT 191.800 145.800 192.200 146.600 ;
        RECT 1.400 140.800 1.800 145.100 ;
        RECT 4.200 140.800 4.600 143.100 ;
        RECT 5.800 140.800 6.200 143.100 ;
        RECT 8.600 140.800 9.000 145.000 ;
        RECT 10.200 140.800 10.600 145.100 ;
        RECT 13.400 140.800 13.800 144.900 ;
        RECT 16.000 140.800 16.400 145.100 ;
        RECT 18.200 140.800 18.600 145.100 ;
        RECT 21.000 140.800 21.400 143.100 ;
        RECT 22.600 140.800 23.000 143.100 ;
        RECT 25.400 140.800 25.800 145.000 ;
        RECT 27.800 140.800 28.200 145.100 ;
        RECT 30.600 140.800 31.000 143.100 ;
        RECT 32.200 140.800 32.600 143.100 ;
        RECT 35.000 140.800 35.400 145.000 ;
        RECT 36.900 140.800 37.300 143.100 ;
        RECT 39.000 140.800 39.400 145.100 ;
        RECT 41.400 140.800 41.800 144.500 ;
        RECT 43.000 140.800 43.400 145.100 ;
        RECT 47.000 140.800 47.500 144.400 ;
        RECT 50.100 141.100 50.600 144.400 ;
        RECT 50.100 140.800 50.500 141.100 ;
        RECT 52.600 140.800 53.000 144.500 ;
        RECT 55.300 140.800 55.700 143.100 ;
        RECT 57.400 140.800 57.800 145.100 ;
        RECT 58.200 140.800 58.600 145.100 ;
        RECT 60.600 140.800 61.000 144.500 ;
        RECT 63.800 140.800 64.200 144.900 ;
        RECT 66.400 140.800 66.800 145.100 ;
        RECT 67.800 140.800 68.200 145.100 ;
        RECT 69.400 140.800 69.800 144.500 ;
        RECT 71.300 140.800 71.700 143.100 ;
        RECT 73.400 140.800 73.800 145.100 ;
        RECT 75.000 140.800 75.400 145.100 ;
        RECT 77.800 140.800 78.200 143.100 ;
        RECT 79.400 140.800 79.800 143.100 ;
        RECT 82.200 140.800 82.600 145.000 ;
        RECT 83.800 140.800 84.200 145.100 ;
        RECT 87.000 140.800 87.400 144.500 ;
        RECT 89.700 140.800 90.100 143.100 ;
        RECT 91.800 140.800 92.200 145.100 ;
        RECT 93.200 140.800 93.600 145.100 ;
        RECT 95.800 140.800 96.200 144.900 ;
        RECT 99.800 140.800 100.200 144.900 ;
        RECT 102.400 140.800 102.800 145.100 ;
        RECT 104.600 140.800 105.000 145.100 ;
        RECT 107.400 140.800 107.800 143.100 ;
        RECT 109.000 140.800 109.400 143.100 ;
        RECT 111.800 140.800 112.200 145.000 ;
        RECT 114.200 140.800 114.600 145.100 ;
        RECT 117.000 140.800 117.400 143.100 ;
        RECT 118.600 140.800 119.000 143.100 ;
        RECT 121.400 140.800 121.800 145.000 ;
        RECT 124.600 140.800 125.000 145.100 ;
        RECT 125.400 140.800 125.800 145.100 ;
        RECT 127.000 140.800 127.400 145.100 ;
        RECT 128.600 140.800 129.000 145.100 ;
        RECT 130.200 140.800 130.600 145.100 ;
        RECT 131.800 140.800 132.200 145.100 ;
        RECT 133.400 140.800 133.800 145.100 ;
        RECT 136.200 140.800 136.600 143.100 ;
        RECT 137.800 140.800 138.200 143.100 ;
        RECT 140.600 140.800 141.000 145.000 ;
        RECT 142.200 140.800 142.600 145.100 ;
        RECT 143.800 140.800 144.200 145.100 ;
        RECT 145.400 140.800 145.800 145.100 ;
        RECT 147.000 140.800 147.400 145.100 ;
        RECT 148.600 140.800 149.000 145.100 ;
        RECT 151.800 140.800 152.200 145.000 ;
        RECT 154.600 140.800 155.000 143.100 ;
        RECT 156.200 140.800 156.600 143.100 ;
        RECT 159.000 140.800 159.400 145.100 ;
        RECT 160.600 140.800 161.000 143.100 ;
        RECT 162.200 140.800 162.600 143.100 ;
        RECT 163.800 140.800 164.200 144.900 ;
        RECT 166.400 140.800 166.800 145.100 ;
        RECT 169.400 140.800 169.800 145.100 ;
        RECT 171.800 140.800 172.200 145.100 ;
        RECT 173.400 140.800 173.800 145.000 ;
        RECT 176.200 140.800 176.600 143.100 ;
        RECT 177.800 140.800 178.200 143.100 ;
        RECT 180.600 140.800 181.000 145.100 ;
        RECT 183.000 140.800 183.400 145.000 ;
        RECT 185.800 140.800 186.200 143.100 ;
        RECT 187.400 140.800 187.800 143.100 ;
        RECT 190.200 140.800 190.600 145.100 ;
        RECT 192.600 140.800 193.000 144.500 ;
        RECT 0.200 140.200 195.800 140.800 ;
        RECT 1.400 135.900 1.800 140.200 ;
        RECT 4.200 137.900 4.600 140.200 ;
        RECT 5.800 137.900 6.200 140.200 ;
        RECT 8.600 136.000 9.000 140.200 ;
        RECT 11.000 136.000 11.400 140.200 ;
        RECT 13.800 137.900 14.200 140.200 ;
        RECT 15.400 137.900 15.800 140.200 ;
        RECT 18.200 135.900 18.600 140.200 ;
        RECT 19.800 135.900 20.200 140.200 ;
        RECT 23.000 136.100 23.400 140.200 ;
        RECT 25.600 135.900 26.000 140.200 ;
        RECT 27.800 136.500 28.200 140.200 ;
        RECT 31.000 135.900 31.400 140.200 ;
        RECT 32.400 135.900 32.800 140.200 ;
        RECT 35.000 136.100 35.400 140.200 ;
        RECT 36.900 137.900 37.300 140.200 ;
        RECT 39.000 135.900 39.400 140.200 ;
        RECT 41.400 136.500 41.800 140.200 ;
        RECT 43.000 137.900 43.400 140.200 ;
        RECT 44.600 138.100 45.000 140.200 ;
        RECT 48.600 136.600 49.100 140.200 ;
        RECT 51.700 139.900 52.100 140.200 ;
        RECT 51.700 136.600 52.200 139.900 ;
        RECT 53.400 135.900 53.800 140.200 ;
        RECT 55.000 136.500 55.400 140.200 ;
        RECT 56.600 135.900 57.000 140.200 ;
        RECT 58.700 137.900 59.100 140.200 ;
        RECT 60.100 137.900 60.500 140.200 ;
        RECT 62.200 135.900 62.600 140.200 ;
        RECT 63.000 137.900 63.400 140.200 ;
        RECT 64.600 138.100 65.000 140.200 ;
        RECT 66.200 137.900 66.600 140.200 ;
        RECT 67.800 138.100 68.200 140.200 ;
        RECT 69.400 137.900 69.800 140.200 ;
        RECT 71.000 137.900 71.400 140.200 ;
        RECT 71.800 137.900 72.200 140.200 ;
        RECT 73.400 138.100 73.800 140.200 ;
        RECT 75.900 139.900 76.300 140.200 ;
        RECT 75.800 136.600 76.300 139.900 ;
        RECT 78.900 136.600 79.400 140.200 ;
        RECT 81.400 136.100 81.800 140.200 ;
        RECT 84.000 135.900 84.400 140.200 ;
        RECT 86.200 136.500 86.600 140.200 ;
        RECT 88.900 137.900 89.300 140.200 ;
        RECT 91.000 135.900 91.400 140.200 ;
        RECT 92.400 135.900 92.800 140.200 ;
        RECT 95.000 136.100 95.400 140.200 ;
        RECT 98.200 135.900 98.600 140.200 ;
        RECT 99.800 136.500 100.200 140.200 ;
        RECT 102.200 136.100 102.600 140.200 ;
        RECT 104.800 135.900 105.200 140.200 ;
        RECT 106.800 135.900 107.200 140.200 ;
        RECT 109.400 136.100 109.800 140.200 ;
        RECT 111.000 137.900 111.400 140.200 ;
        RECT 113.200 135.900 113.600 140.200 ;
        RECT 115.800 136.100 116.200 140.200 ;
        RECT 118.200 136.100 118.600 140.200 ;
        RECT 120.800 135.900 121.200 140.200 ;
        RECT 122.800 135.900 123.200 140.200 ;
        RECT 125.400 136.100 125.800 140.200 ;
        RECT 127.800 136.100 128.200 140.200 ;
        RECT 130.400 135.900 130.800 140.200 ;
        RECT 133.400 136.500 133.800 140.200 ;
        RECT 135.000 135.900 135.400 140.200 ;
        RECT 137.100 137.900 137.500 140.200 ;
        RECT 139.300 135.900 139.700 140.200 ;
        RECT 141.400 137.900 141.800 140.200 ;
        RECT 143.000 137.900 143.400 140.200 ;
        RECT 143.800 137.900 144.200 140.200 ;
        RECT 145.400 137.900 145.800 140.200 ;
        RECT 146.500 137.900 146.900 140.200 ;
        RECT 148.600 135.900 149.000 140.200 ;
        RECT 151.000 137.900 151.400 140.200 ;
        RECT 152.600 135.900 153.000 140.200 ;
        RECT 154.700 137.900 155.100 140.200 ;
        RECT 155.800 135.900 156.200 140.200 ;
        RECT 158.200 136.500 158.600 140.200 ;
        RECT 160.600 135.900 161.000 140.200 ;
        RECT 162.700 137.900 163.100 140.200 ;
        RECT 164.100 137.900 164.500 140.200 ;
        RECT 166.200 135.900 166.600 140.200 ;
        RECT 168.600 136.500 169.000 140.200 ;
        RECT 171.000 136.000 171.400 140.200 ;
        RECT 173.800 137.900 174.200 140.200 ;
        RECT 175.400 137.900 175.800 140.200 ;
        RECT 178.200 135.900 178.600 140.200 ;
        RECT 180.600 135.900 181.000 140.200 ;
        RECT 183.400 137.900 183.800 140.200 ;
        RECT 185.000 137.900 185.400 140.200 ;
        RECT 187.800 136.000 188.200 140.200 ;
        RECT 190.200 136.500 190.600 140.200 ;
        RECT 192.600 136.500 193.000 140.200 ;
        RECT 1.400 120.800 1.800 125.100 ;
        RECT 4.200 120.800 4.600 123.100 ;
        RECT 5.800 120.800 6.200 123.100 ;
        RECT 8.600 120.800 9.000 125.000 ;
        RECT 11.000 120.800 11.400 125.100 ;
        RECT 13.800 120.800 14.200 123.100 ;
        RECT 15.400 120.800 15.800 123.100 ;
        RECT 18.200 120.800 18.600 125.000 ;
        RECT 20.600 120.800 21.000 125.000 ;
        RECT 23.400 120.800 23.800 123.100 ;
        RECT 25.000 120.800 25.400 123.100 ;
        RECT 27.800 120.800 28.200 125.100 ;
        RECT 29.400 120.800 29.800 125.100 ;
        RECT 31.000 120.800 31.400 123.100 ;
        RECT 32.600 120.800 33.000 123.100 ;
        RECT 33.400 120.800 33.800 123.100 ;
        RECT 35.300 120.800 35.700 123.100 ;
        RECT 37.400 120.800 37.800 125.100 ;
        RECT 38.200 120.800 38.600 125.100 ;
        RECT 41.400 120.800 41.800 122.900 ;
        RECT 43.000 120.800 43.400 123.100 ;
        RECT 43.800 120.800 44.200 123.100 ;
        RECT 47.300 120.800 47.700 123.100 ;
        RECT 49.400 120.800 49.800 125.100 ;
        RECT 51.800 120.800 52.200 125.100 ;
        RECT 52.600 120.800 53.000 123.100 ;
        RECT 54.200 120.800 54.600 123.100 ;
        RECT 55.800 120.800 56.200 122.900 ;
        RECT 57.400 120.800 57.800 125.100 ;
        RECT 59.800 120.800 60.200 123.100 ;
        RECT 61.400 120.800 61.800 123.100 ;
        RECT 62.200 120.800 62.600 123.100 ;
        RECT 63.800 120.800 64.200 123.100 ;
        RECT 65.400 120.800 65.800 122.900 ;
        RECT 67.000 120.800 67.400 123.100 ;
        RECT 69.400 120.800 69.800 125.100 ;
        RECT 71.000 120.800 71.400 124.100 ;
        RECT 76.600 120.800 77.000 125.100 ;
        RECT 79.000 120.800 79.400 125.100 ;
        RECT 81.100 120.800 81.500 123.100 ;
        RECT 82.200 120.800 82.600 123.100 ;
        RECT 83.800 120.800 84.200 123.100 ;
        RECT 84.600 120.800 85.000 125.100 ;
        RECT 86.200 120.800 86.600 125.100 ;
        RECT 87.000 120.800 87.400 125.100 ;
        RECT 90.200 120.800 90.600 123.100 ;
        RECT 91.800 120.800 92.200 125.100 ;
        RECT 94.600 120.800 95.000 123.100 ;
        RECT 96.200 120.800 96.600 123.100 ;
        RECT 99.000 120.800 99.400 125.000 ;
        RECT 102.200 120.800 102.600 125.100 ;
        RECT 103.800 120.800 104.200 125.100 ;
        RECT 105.400 120.800 105.800 125.100 ;
        RECT 107.000 120.800 107.400 125.100 ;
        RECT 108.600 120.800 109.000 125.100 ;
        RECT 109.400 120.800 109.800 125.100 ;
        RECT 111.000 120.800 111.400 124.500 ;
        RECT 113.400 120.800 113.800 124.900 ;
        RECT 116.000 120.800 116.400 125.100 ;
        RECT 117.400 120.800 117.800 123.100 ;
        RECT 119.000 120.800 119.400 125.100 ;
        RECT 120.600 120.800 121.000 124.500 ;
        RECT 122.200 120.800 122.600 125.100 ;
        RECT 123.800 120.800 124.200 125.100 ;
        RECT 125.400 120.800 125.800 125.100 ;
        RECT 127.000 120.800 127.400 125.100 ;
        RECT 128.600 120.800 129.000 125.100 ;
        RECT 130.200 120.800 130.600 124.500 ;
        RECT 131.800 120.800 132.200 125.100 ;
        RECT 133.400 120.800 133.800 124.500 ;
        RECT 135.000 120.800 135.400 125.100 ;
        RECT 136.600 120.800 137.000 125.100 ;
        RECT 137.400 120.800 137.800 125.100 ;
        RECT 139.500 120.800 139.900 123.100 ;
        RECT 142.200 120.800 142.600 124.500 ;
        RECT 143.800 120.800 144.200 123.100 ;
        RECT 145.400 120.800 145.800 123.100 ;
        RECT 146.200 120.800 146.600 125.100 ;
        RECT 151.800 120.800 152.200 125.100 ;
        RECT 153.400 120.800 153.800 124.500 ;
        RECT 156.600 120.800 157.000 122.900 ;
        RECT 158.200 120.800 158.600 123.100 ;
        RECT 159.000 120.800 159.400 123.100 ;
        RECT 160.600 120.800 161.000 123.100 ;
        RECT 163.000 120.800 163.400 125.100 ;
        RECT 164.100 120.800 164.500 123.100 ;
        RECT 166.200 120.800 166.600 125.100 ;
        RECT 167.800 120.800 168.300 124.400 ;
        RECT 170.900 121.100 171.400 124.400 ;
        RECT 170.900 120.800 171.300 121.100 ;
        RECT 173.400 120.800 173.800 125.100 ;
        RECT 176.200 120.800 176.600 123.100 ;
        RECT 177.800 120.800 178.200 123.100 ;
        RECT 180.600 120.800 181.000 125.000 ;
        RECT 182.800 120.800 183.200 125.100 ;
        RECT 185.400 120.800 185.800 124.900 ;
        RECT 187.000 120.800 187.400 123.100 ;
        RECT 188.600 120.800 189.000 125.100 ;
        RECT 191.800 120.800 192.200 124.500 ;
        RECT 193.400 120.800 193.800 125.100 ;
        RECT 0.200 120.200 195.800 120.800 ;
        RECT 1.400 115.900 1.800 120.200 ;
        RECT 4.200 117.900 4.600 120.200 ;
        RECT 5.800 117.900 6.200 120.200 ;
        RECT 8.600 116.000 9.000 120.200 ;
        RECT 10.200 115.900 10.600 120.200 ;
        RECT 12.600 117.900 13.000 120.200 ;
        RECT 14.200 116.100 14.600 120.200 ;
        RECT 16.600 116.000 17.000 120.200 ;
        RECT 19.400 117.900 19.800 120.200 ;
        RECT 21.000 117.900 21.400 120.200 ;
        RECT 23.800 115.900 24.200 120.200 ;
        RECT 26.200 115.900 26.600 120.200 ;
        RECT 29.000 117.900 29.400 120.200 ;
        RECT 30.600 117.900 31.000 120.200 ;
        RECT 33.400 116.000 33.800 120.200 ;
        RECT 35.000 115.900 35.400 120.200 ;
        RECT 37.100 117.900 37.500 120.200 ;
        RECT 39.800 116.500 40.200 120.200 ;
        RECT 41.400 115.900 41.800 120.200 ;
        RECT 44.600 118.100 45.000 120.200 ;
        RECT 46.200 117.900 46.600 120.200 ;
        RECT 49.400 118.100 49.800 120.200 ;
        RECT 51.000 117.900 51.400 120.200 ;
        RECT 52.600 118.100 53.000 120.200 ;
        RECT 54.200 117.900 54.600 120.200 ;
        RECT 55.800 117.900 56.200 120.200 ;
        RECT 56.600 117.900 57.000 120.200 ;
        RECT 58.200 117.900 58.600 120.200 ;
        RECT 59.300 117.900 59.700 120.200 ;
        RECT 61.400 115.900 61.800 120.200 ;
        RECT 63.000 117.900 63.400 120.200 ;
        RECT 64.600 116.100 65.000 120.200 ;
        RECT 66.200 117.900 66.600 120.200 ;
        RECT 67.000 115.900 67.400 120.200 ;
        RECT 70.200 115.900 70.600 120.200 ;
        RECT 73.000 117.900 73.400 120.200 ;
        RECT 74.600 117.900 75.000 120.200 ;
        RECT 77.400 116.000 77.800 120.200 ;
        RECT 79.800 117.900 80.200 120.200 ;
        RECT 80.600 115.900 81.000 120.200 ;
        RECT 82.700 117.900 83.100 120.200 ;
        RECT 83.800 117.900 84.200 120.200 ;
        RECT 85.400 117.900 85.800 120.200 ;
        RECT 87.000 116.100 87.400 120.200 ;
        RECT 89.600 115.900 90.000 120.200 ;
        RECT 92.600 115.900 93.000 120.200 ;
        RECT 95.800 115.900 96.200 120.200 ;
        RECT 98.600 117.900 99.000 120.200 ;
        RECT 100.200 117.900 100.600 120.200 ;
        RECT 103.000 116.000 103.400 120.200 ;
        RECT 105.400 116.000 105.800 120.200 ;
        RECT 108.200 117.900 108.600 120.200 ;
        RECT 109.800 117.900 110.200 120.200 ;
        RECT 112.600 115.900 113.000 120.200 ;
        RECT 115.000 115.900 115.400 120.200 ;
        RECT 117.800 117.900 118.200 120.200 ;
        RECT 119.400 117.900 119.800 120.200 ;
        RECT 122.200 116.000 122.600 120.200 ;
        RECT 123.800 115.900 124.200 120.200 ;
        RECT 126.800 115.900 127.200 120.200 ;
        RECT 129.400 116.100 129.800 120.200 ;
        RECT 131.000 117.900 131.400 120.200 ;
        RECT 132.600 117.900 133.000 120.200 ;
        RECT 133.400 115.900 133.800 120.200 ;
        RECT 135.800 117.900 136.200 120.200 ;
        RECT 137.400 117.900 137.800 120.200 ;
        RECT 138.500 117.900 138.900 120.200 ;
        RECT 140.600 115.900 141.000 120.200 ;
        RECT 142.200 117.900 142.600 120.200 ;
        RECT 143.800 117.900 144.200 120.200 ;
        RECT 147.000 115.900 147.400 120.200 ;
        RECT 149.800 117.900 150.200 120.200 ;
        RECT 151.400 117.900 151.800 120.200 ;
        RECT 154.200 116.000 154.600 120.200 ;
        RECT 155.800 117.900 156.200 120.200 ;
        RECT 157.400 116.100 157.800 120.200 ;
        RECT 159.800 115.900 160.200 120.200 ;
        RECT 162.600 117.900 163.000 120.200 ;
        RECT 164.200 117.900 164.600 120.200 ;
        RECT 167.000 116.000 167.400 120.200 ;
        RECT 169.400 115.900 169.800 120.200 ;
        RECT 172.200 117.900 172.600 120.200 ;
        RECT 173.800 117.900 174.200 120.200 ;
        RECT 176.600 116.000 177.000 120.200 ;
        RECT 178.800 115.900 179.200 120.200 ;
        RECT 181.400 116.100 181.800 120.200 ;
        RECT 183.300 117.900 183.700 120.200 ;
        RECT 185.400 115.900 185.800 120.200 ;
        RECT 187.000 116.500 187.400 120.200 ;
        RECT 189.400 116.500 189.800 120.200 ;
        RECT 192.600 116.500 193.000 120.200 ;
        RECT 0.600 100.800 1.000 103.100 ;
        RECT 2.200 100.800 2.600 103.100 ;
        RECT 3.300 100.800 3.700 103.100 ;
        RECT 5.400 100.800 5.800 105.100 ;
        RECT 7.000 100.800 7.400 103.100 ;
        RECT 7.800 100.800 8.200 103.100 ;
        RECT 9.400 100.800 9.800 104.900 ;
        RECT 11.000 100.800 11.400 105.100 ;
        RECT 13.400 100.800 13.800 105.100 ;
        RECT 16.600 100.800 17.000 105.100 ;
        RECT 17.400 100.800 17.800 103.100 ;
        RECT 19.000 100.800 19.400 103.100 ;
        RECT 20.100 100.800 20.500 103.100 ;
        RECT 22.200 100.800 22.600 105.100 ;
        RECT 23.800 100.800 24.200 103.100 ;
        RECT 25.400 101.100 25.900 104.400 ;
        RECT 25.500 100.800 25.900 101.100 ;
        RECT 28.500 100.800 29.000 104.400 ;
        RECT 30.200 100.800 30.600 103.100 ;
        RECT 31.800 100.800 32.200 103.100 ;
        RECT 32.900 100.800 33.300 103.100 ;
        RECT 35.000 100.800 35.400 105.100 ;
        RECT 36.600 100.800 37.000 103.100 ;
        RECT 37.400 100.800 37.800 103.100 ;
        RECT 39.000 100.800 39.400 103.100 ;
        RECT 39.800 100.800 40.200 103.100 ;
        RECT 41.400 100.800 41.800 102.900 ;
        RECT 45.400 100.800 45.800 104.100 ;
        RECT 51.000 100.800 51.400 105.100 ;
        RECT 52.600 100.800 53.000 104.500 ;
        RECT 55.000 100.800 55.400 104.900 ;
        RECT 57.600 100.800 58.000 105.100 ;
        RECT 59.000 100.800 59.400 103.100 ;
        RECT 60.600 100.800 61.000 103.100 ;
        RECT 61.400 100.800 61.800 105.100 ;
        RECT 64.600 100.800 65.000 105.100 ;
        RECT 65.400 100.800 65.800 105.100 ;
        RECT 67.800 100.800 68.200 103.100 ;
        RECT 69.400 100.800 69.800 104.900 ;
        RECT 71.300 100.800 71.700 103.100 ;
        RECT 73.400 100.800 73.800 105.100 ;
        RECT 75.000 100.800 75.400 103.100 ;
        RECT 75.800 100.800 76.200 105.100 ;
        RECT 77.400 100.800 77.800 105.100 ;
        RECT 79.000 100.800 79.400 105.100 ;
        RECT 80.600 100.800 81.000 105.100 ;
        RECT 82.200 100.800 82.600 105.100 ;
        RECT 83.800 100.800 84.200 105.100 ;
        RECT 86.600 100.800 87.000 103.100 ;
        RECT 88.200 100.800 88.600 103.100 ;
        RECT 91.000 100.800 91.400 105.000 ;
        RECT 95.000 100.800 95.400 105.100 ;
        RECT 97.800 100.800 98.200 103.100 ;
        RECT 99.400 100.800 99.800 103.100 ;
        RECT 102.200 100.800 102.600 105.000 ;
        RECT 104.600 100.800 105.000 105.100 ;
        RECT 107.400 100.800 107.800 103.100 ;
        RECT 109.000 100.800 109.400 103.100 ;
        RECT 111.800 100.800 112.200 105.000 ;
        RECT 113.400 100.800 113.800 105.100 ;
        RECT 115.800 100.800 116.200 105.100 ;
        RECT 117.400 100.800 117.800 105.100 ;
        RECT 119.000 100.800 119.400 105.100 ;
        RECT 120.600 100.800 121.000 105.100 ;
        RECT 122.200 100.800 122.600 105.100 ;
        RECT 123.800 100.800 124.200 104.900 ;
        RECT 126.400 100.800 126.800 105.100 ;
        RECT 128.600 100.800 129.000 105.000 ;
        RECT 131.400 100.800 131.800 103.100 ;
        RECT 133.000 100.800 133.400 103.100 ;
        RECT 135.800 100.800 136.200 105.100 ;
        RECT 138.200 100.800 138.600 105.000 ;
        RECT 141.000 100.800 141.400 103.100 ;
        RECT 142.600 100.800 143.000 103.100 ;
        RECT 145.400 100.800 145.800 105.100 ;
        RECT 147.000 100.800 147.400 103.100 ;
        RECT 148.600 100.800 149.000 103.100 ;
        RECT 151.300 100.800 151.700 103.100 ;
        RECT 153.400 100.800 153.800 105.100 ;
        RECT 155.000 100.800 155.400 103.100 ;
        RECT 155.800 100.800 156.200 105.100 ;
        RECT 158.200 100.800 158.600 105.100 ;
        RECT 161.400 100.800 161.800 105.100 ;
        RECT 162.200 100.800 162.600 105.100 ;
        RECT 165.400 100.800 165.800 104.900 ;
        RECT 167.000 100.800 167.400 103.100 ;
        RECT 168.600 100.800 169.000 104.900 ;
        RECT 171.200 100.800 171.600 105.100 ;
        RECT 174.200 100.800 174.600 105.100 ;
        RECT 175.000 100.800 175.400 105.100 ;
        RECT 176.600 100.800 177.000 105.100 ;
        RECT 178.200 100.800 178.600 105.100 ;
        RECT 179.800 100.800 180.200 105.100 ;
        RECT 181.400 100.800 181.800 105.100 ;
        RECT 182.800 100.800 183.200 105.100 ;
        RECT 185.400 100.800 185.800 104.900 ;
        RECT 187.800 100.800 188.200 104.900 ;
        RECT 190.400 100.800 190.800 105.100 ;
        RECT 193.100 100.800 193.500 105.100 ;
        RECT 0.200 100.200 195.800 100.800 ;
        RECT 1.400 96.500 1.800 100.200 ;
        RECT 3.300 97.900 3.700 100.200 ;
        RECT 5.400 95.900 5.800 100.200 ;
        RECT 7.000 97.900 7.400 100.200 ;
        RECT 8.700 99.900 9.100 100.200 ;
        RECT 8.600 96.600 9.100 99.900 ;
        RECT 11.700 96.600 12.200 100.200 ;
        RECT 14.200 95.900 14.600 100.200 ;
        RECT 17.000 97.900 17.400 100.200 ;
        RECT 18.600 97.900 19.000 100.200 ;
        RECT 21.400 96.000 21.800 100.200 ;
        RECT 27.800 96.900 28.200 100.200 ;
        RECT 31.000 96.500 31.400 100.200 ;
        RECT 32.600 95.900 33.000 100.200 ;
        RECT 34.700 97.900 35.100 100.200 ;
        RECT 35.800 95.900 36.200 100.200 ;
        RECT 37.900 97.900 38.300 100.200 ;
        RECT 40.600 95.900 41.000 100.200 ;
        RECT 41.400 97.900 41.800 100.200 ;
        RECT 43.000 97.900 43.400 100.200 ;
        RECT 45.400 96.500 45.800 100.200 ;
        RECT 49.400 96.600 49.900 100.200 ;
        RECT 52.500 99.900 52.900 100.200 ;
        RECT 52.500 96.600 53.000 99.900 ;
        RECT 54.200 97.900 54.600 100.200 ;
        RECT 55.800 97.900 56.200 100.200 ;
        RECT 57.400 96.900 57.800 100.200 ;
        RECT 63.800 96.600 64.300 100.200 ;
        RECT 66.900 99.900 67.300 100.200 ;
        RECT 66.900 96.600 67.400 99.900 ;
        RECT 68.600 97.900 69.000 100.200 ;
        RECT 70.200 95.900 70.600 100.200 ;
        RECT 72.300 97.900 72.700 100.200 ;
        RECT 74.200 96.100 74.600 100.200 ;
        RECT 76.800 95.900 77.200 100.200 ;
        RECT 79.800 95.900 80.200 100.200 ;
        RECT 81.400 96.100 81.800 100.200 ;
        RECT 84.000 95.900 84.400 100.200 ;
        RECT 87.000 95.900 87.400 100.200 ;
        RECT 88.600 95.900 89.000 100.200 ;
        RECT 91.400 97.900 91.800 100.200 ;
        RECT 93.000 97.900 93.400 100.200 ;
        RECT 95.800 96.000 96.200 100.200 ;
        RECT 99.000 95.900 99.400 100.200 ;
        RECT 100.600 95.900 101.000 100.200 ;
        RECT 102.200 95.900 102.600 100.200 ;
        RECT 103.800 95.900 104.200 100.200 ;
        RECT 105.400 95.900 105.800 100.200 ;
        RECT 106.200 95.900 106.600 100.200 ;
        RECT 109.400 96.100 109.800 100.200 ;
        RECT 112.000 95.900 112.400 100.200 ;
        RECT 113.700 97.900 114.100 100.200 ;
        RECT 115.800 95.900 116.200 100.200 ;
        RECT 116.600 97.900 117.000 100.200 ;
        RECT 118.200 97.900 118.600 100.200 ;
        RECT 119.800 97.900 120.200 100.200 ;
        RECT 120.900 97.900 121.300 100.200 ;
        RECT 123.000 95.900 123.400 100.200 ;
        RECT 124.600 97.900 125.000 100.200 ;
        RECT 126.200 96.600 126.700 100.200 ;
        RECT 129.300 99.900 129.700 100.200 ;
        RECT 129.300 96.600 129.800 99.900 ;
        RECT 131.800 96.900 132.200 100.200 ;
        RECT 138.300 99.900 138.700 100.200 ;
        RECT 138.200 96.600 138.700 99.900 ;
        RECT 141.300 96.600 141.800 100.200 ;
        RECT 143.800 95.900 144.200 100.200 ;
        RECT 146.600 97.900 147.000 100.200 ;
        RECT 148.200 97.900 148.600 100.200 ;
        RECT 151.000 96.000 151.400 100.200 ;
        RECT 155.000 95.900 155.400 100.200 ;
        RECT 157.800 97.900 158.200 100.200 ;
        RECT 159.400 97.900 159.800 100.200 ;
        RECT 162.200 96.000 162.600 100.200 ;
        RECT 164.600 96.000 165.000 100.200 ;
        RECT 167.400 97.900 167.800 100.200 ;
        RECT 169.000 97.900 169.400 100.200 ;
        RECT 171.800 95.900 172.200 100.200 ;
        RECT 174.200 95.900 174.600 100.200 ;
        RECT 177.000 97.900 177.400 100.200 ;
        RECT 178.600 97.900 179.000 100.200 ;
        RECT 181.400 96.000 181.800 100.200 ;
        RECT 183.800 96.000 184.200 100.200 ;
        RECT 186.600 97.900 187.000 100.200 ;
        RECT 188.200 97.900 188.600 100.200 ;
        RECT 191.000 95.900 191.400 100.200 ;
        RECT 193.400 96.500 193.800 100.200 ;
        RECT 188.600 85.800 189.000 86.600 ;
        RECT 0.600 80.800 1.000 83.100 ;
        RECT 2.200 80.800 2.600 83.100 ;
        RECT 3.600 80.800 4.000 85.100 ;
        RECT 6.200 80.800 6.600 84.900 ;
        RECT 8.600 80.800 9.000 84.900 ;
        RECT 11.200 80.800 11.600 85.100 ;
        RECT 13.400 80.800 13.800 85.100 ;
        RECT 16.200 80.800 16.600 83.100 ;
        RECT 17.800 80.800 18.200 83.100 ;
        RECT 20.600 80.800 21.000 85.000 ;
        RECT 22.200 80.800 22.600 85.100 ;
        RECT 23.800 80.800 24.200 84.500 ;
        RECT 26.200 80.800 26.600 84.500 ;
        RECT 27.800 80.800 28.200 85.100 ;
        RECT 28.600 80.800 29.000 85.100 ;
        RECT 31.800 80.800 32.200 85.100 ;
        RECT 32.600 80.800 33.000 83.100 ;
        RECT 34.200 80.800 34.600 83.100 ;
        RECT 35.000 80.800 35.400 83.100 ;
        RECT 36.600 80.800 37.000 83.100 ;
        RECT 38.200 80.800 38.600 83.100 ;
        RECT 39.000 80.800 39.400 83.100 ;
        RECT 40.600 80.800 41.000 83.100 ;
        RECT 41.700 80.800 42.100 83.100 ;
        RECT 43.800 80.800 44.200 85.100 ;
        RECT 44.600 80.800 45.000 85.100 ;
        RECT 49.400 81.100 49.900 84.400 ;
        RECT 49.500 80.800 49.900 81.100 ;
        RECT 52.500 80.800 53.000 84.400 ;
        RECT 54.500 80.800 54.900 83.100 ;
        RECT 56.600 80.800 57.000 85.100 ;
        RECT 58.200 80.800 58.600 83.100 ;
        RECT 59.000 80.800 59.400 83.100 ;
        RECT 60.600 80.800 61.000 82.900 ;
        RECT 63.000 80.800 63.400 85.100 ;
        RECT 65.800 80.800 66.200 83.100 ;
        RECT 67.400 80.800 67.800 83.100 ;
        RECT 70.200 80.800 70.600 85.000 ;
        RECT 71.800 80.800 72.200 83.100 ;
        RECT 73.400 80.800 73.800 83.100 ;
        RECT 75.000 80.800 75.400 85.100 ;
        RECT 77.800 80.800 78.200 83.100 ;
        RECT 79.400 80.800 79.800 83.100 ;
        RECT 82.200 80.800 82.600 85.000 ;
        RECT 83.800 80.800 84.200 85.100 ;
        RECT 85.400 80.800 85.800 84.500 ;
        RECT 87.800 80.800 88.200 85.100 ;
        RECT 90.600 80.800 91.000 83.100 ;
        RECT 92.200 80.800 92.600 83.100 ;
        RECT 95.000 80.800 95.400 85.000 ;
        RECT 99.000 80.800 99.400 85.100 ;
        RECT 101.800 80.800 102.200 83.100 ;
        RECT 103.400 80.800 103.800 83.100 ;
        RECT 106.200 80.800 106.600 85.000 ;
        RECT 108.600 80.800 109.000 85.100 ;
        RECT 111.400 80.800 111.800 83.100 ;
        RECT 113.000 80.800 113.400 83.100 ;
        RECT 115.800 80.800 116.200 85.000 ;
        RECT 117.400 80.800 117.800 85.100 ;
        RECT 119.800 80.800 120.200 83.100 ;
        RECT 121.400 80.800 121.800 83.100 ;
        RECT 123.000 80.800 123.400 84.900 ;
        RECT 125.600 80.800 126.000 85.100 ;
        RECT 127.800 80.800 128.200 85.100 ;
        RECT 130.600 80.800 131.000 83.100 ;
        RECT 132.200 80.800 132.600 83.100 ;
        RECT 135.000 80.800 135.400 85.000 ;
        RECT 136.600 80.800 137.000 85.100 ;
        RECT 139.600 80.800 140.000 85.100 ;
        RECT 142.200 80.800 142.600 84.900 ;
        RECT 146.200 80.800 146.600 85.100 ;
        RECT 149.000 80.800 149.400 83.100 ;
        RECT 150.600 80.800 151.000 83.100 ;
        RECT 153.400 80.800 153.800 85.000 ;
        RECT 155.800 80.800 156.200 84.500 ;
        RECT 157.400 80.800 157.800 85.100 ;
        RECT 159.500 80.800 159.900 83.100 ;
        RECT 160.600 80.800 161.000 83.100 ;
        RECT 162.200 80.800 162.600 83.100 ;
        RECT 163.800 80.800 164.200 82.900 ;
        RECT 165.400 80.800 165.800 83.100 ;
        RECT 166.200 80.800 166.600 83.100 ;
        RECT 167.800 80.800 168.200 82.900 ;
        RECT 169.400 80.800 169.800 85.100 ;
        RECT 171.800 80.800 172.200 85.100 ;
        RECT 173.400 80.800 173.800 85.100 ;
        RECT 175.500 80.800 175.900 83.100 ;
        RECT 176.600 80.800 177.000 85.100 ;
        RECT 180.600 80.800 181.000 85.100 ;
        RECT 182.200 80.800 182.700 84.400 ;
        RECT 185.300 81.100 185.800 84.400 ;
        RECT 185.300 80.800 185.700 81.100 ;
        RECT 187.800 80.800 188.200 84.500 ;
        RECT 190.200 80.800 190.600 84.500 ;
        RECT 192.600 80.800 193.000 84.500 ;
        RECT 0.200 80.200 195.800 80.800 ;
        RECT 0.600 75.900 1.000 80.200 ;
        RECT 2.200 75.900 2.600 80.200 ;
        RECT 3.800 75.900 4.200 80.200 ;
        RECT 5.400 75.900 5.800 80.200 ;
        RECT 7.000 75.900 7.400 80.200 ;
        RECT 9.400 75.900 9.800 80.200 ;
        RECT 11.000 75.900 11.400 80.200 ;
        RECT 13.800 77.900 14.200 80.200 ;
        RECT 15.400 77.900 15.800 80.200 ;
        RECT 18.200 76.000 18.600 80.200 ;
        RECT 20.600 76.000 21.000 80.200 ;
        RECT 23.400 77.900 23.800 80.200 ;
        RECT 25.000 77.900 25.400 80.200 ;
        RECT 27.800 75.900 28.200 80.200 ;
        RECT 29.400 75.900 29.800 80.200 ;
        RECT 32.600 75.900 33.000 80.200 ;
        RECT 35.400 77.900 35.800 80.200 ;
        RECT 37.000 77.900 37.400 80.200 ;
        RECT 39.800 76.000 40.200 80.200 ;
        RECT 41.400 75.900 41.800 80.200 ;
        RECT 43.800 77.900 44.200 80.200 ;
        RECT 45.400 77.900 45.800 80.200 ;
        RECT 49.400 75.900 49.800 80.200 ;
        RECT 51.000 77.900 51.400 80.200 ;
        RECT 51.800 77.900 52.200 80.200 ;
        RECT 53.400 77.900 53.800 80.200 ;
        RECT 54.500 77.900 54.900 80.200 ;
        RECT 56.600 75.900 57.000 80.200 ;
        RECT 58.700 75.900 59.100 80.200 ;
        RECT 61.400 76.500 61.800 80.200 ;
        RECT 64.600 78.100 65.000 80.200 ;
        RECT 66.200 77.900 66.600 80.200 ;
        RECT 67.800 75.900 68.200 80.200 ;
        RECT 70.600 77.900 71.000 80.200 ;
        RECT 72.200 77.900 72.600 80.200 ;
        RECT 75.000 76.000 75.400 80.200 ;
        RECT 77.400 76.500 77.800 80.200 ;
        RECT 79.800 75.900 80.200 80.200 ;
        RECT 81.900 77.900 82.300 80.200 ;
        RECT 83.300 77.900 83.700 80.200 ;
        RECT 85.400 75.900 85.800 80.200 ;
        RECT 86.500 77.900 86.900 80.200 ;
        RECT 88.600 75.900 89.000 80.200 ;
        RECT 89.400 75.900 89.800 80.200 ;
        RECT 91.000 76.500 91.400 80.200 ;
        RECT 93.200 75.900 93.600 80.200 ;
        RECT 95.800 76.100 96.200 80.200 ;
        RECT 99.800 76.500 100.200 80.200 ;
        RECT 101.400 75.900 101.800 80.200 ;
        RECT 102.200 75.900 102.600 80.200 ;
        RECT 103.800 75.900 104.200 80.200 ;
        RECT 105.400 75.900 105.800 80.200 ;
        RECT 107.000 76.000 107.400 80.200 ;
        RECT 109.800 77.900 110.200 80.200 ;
        RECT 111.400 77.900 111.800 80.200 ;
        RECT 114.200 75.900 114.600 80.200 ;
        RECT 116.600 76.000 117.000 80.200 ;
        RECT 119.400 77.900 119.800 80.200 ;
        RECT 121.000 77.900 121.400 80.200 ;
        RECT 123.800 75.900 124.200 80.200 ;
        RECT 127.000 75.900 127.400 80.200 ;
        RECT 127.800 75.900 128.200 80.200 ;
        RECT 129.400 75.900 129.800 80.200 ;
        RECT 131.000 75.900 131.400 80.200 ;
        RECT 132.600 75.900 133.000 80.200 ;
        RECT 134.200 75.900 134.600 80.200 ;
        RECT 135.000 75.900 135.400 80.200 ;
        RECT 136.600 75.900 137.000 80.200 ;
        RECT 138.200 75.900 138.600 80.200 ;
        RECT 139.800 76.000 140.200 80.200 ;
        RECT 142.600 77.900 143.000 80.200 ;
        RECT 144.200 77.900 144.600 80.200 ;
        RECT 147.000 75.900 147.400 80.200 ;
        RECT 151.000 76.500 151.400 80.200 ;
        RECT 152.600 77.900 153.000 80.200 ;
        RECT 155.000 76.000 155.400 80.200 ;
        RECT 157.800 77.900 158.200 80.200 ;
        RECT 159.400 77.900 159.800 80.200 ;
        RECT 162.200 75.900 162.600 80.200 ;
        RECT 165.400 75.900 165.800 80.200 ;
        RECT 166.200 77.900 166.600 80.200 ;
        RECT 167.800 77.900 168.200 80.200 ;
        RECT 168.600 77.900 169.000 80.200 ;
        RECT 170.500 77.900 170.900 80.200 ;
        RECT 172.600 75.900 173.000 80.200 ;
        RECT 173.400 77.900 173.800 80.200 ;
        RECT 176.600 75.900 177.000 80.200 ;
        RECT 179.000 76.500 179.400 80.200 ;
        RECT 180.600 77.900 181.000 80.200 ;
        RECT 182.200 77.900 182.600 80.200 ;
        RECT 183.800 77.900 184.200 80.200 ;
        RECT 185.400 76.000 185.800 80.200 ;
        RECT 188.200 77.900 188.600 80.200 ;
        RECT 189.800 77.900 190.200 80.200 ;
        RECT 192.600 75.900 193.000 80.200 ;
        RECT 150.200 74.400 150.600 75.200 ;
        RECT 189.400 65.800 189.800 66.600 ;
        RECT 191.800 65.800 192.200 66.600 ;
        RECT 1.400 60.800 1.800 64.500 ;
        RECT 3.000 60.800 3.400 65.100 ;
        RECT 4.600 60.800 5.000 65.100 ;
        RECT 6.200 60.800 6.600 65.100 ;
        RECT 7.800 60.800 8.200 65.100 ;
        RECT 9.400 60.800 9.800 65.100 ;
        RECT 11.000 60.800 11.400 65.100 ;
        RECT 13.800 60.800 14.200 63.100 ;
        RECT 15.400 60.800 15.800 63.100 ;
        RECT 18.200 60.800 18.600 65.000 ;
        RECT 20.100 60.800 20.500 63.100 ;
        RECT 22.200 60.800 22.600 65.100 ;
        RECT 23.800 60.800 24.200 63.100 ;
        RECT 25.400 60.800 25.800 65.000 ;
        RECT 28.200 60.800 28.600 63.100 ;
        RECT 29.800 60.800 30.200 63.100 ;
        RECT 32.600 60.800 33.000 65.100 ;
        RECT 34.500 60.800 34.900 63.100 ;
        RECT 36.600 60.800 37.000 65.100 ;
        RECT 38.200 60.800 38.600 63.100 ;
        RECT 39.800 60.800 40.200 65.000 ;
        RECT 42.600 60.800 43.000 63.100 ;
        RECT 44.200 60.800 44.600 63.100 ;
        RECT 47.000 60.800 47.400 65.100 ;
        RECT 50.200 60.800 50.600 63.100 ;
        RECT 51.800 60.800 52.200 63.100 ;
        RECT 53.400 60.800 53.800 63.100 ;
        RECT 55.000 60.800 55.400 64.500 ;
        RECT 57.700 60.800 58.100 63.100 ;
        RECT 59.800 60.800 60.200 65.100 ;
        RECT 62.200 60.800 62.600 65.100 ;
        RECT 63.800 60.800 64.200 65.100 ;
        RECT 66.600 60.800 67.000 63.100 ;
        RECT 68.200 60.800 68.600 63.100 ;
        RECT 71.000 60.800 71.400 65.000 ;
        RECT 73.400 60.800 73.800 64.900 ;
        RECT 76.000 60.800 76.400 65.100 ;
        RECT 78.200 60.800 78.600 65.100 ;
        RECT 81.000 60.800 81.400 63.100 ;
        RECT 82.600 60.800 83.000 63.100 ;
        RECT 85.400 60.800 85.800 65.000 ;
        RECT 87.000 60.800 87.400 65.100 ;
        RECT 90.200 60.800 90.600 65.000 ;
        RECT 93.000 60.800 93.400 63.100 ;
        RECT 94.600 60.800 95.000 63.100 ;
        RECT 97.400 60.800 97.800 65.100 ;
        RECT 101.400 60.800 101.800 65.100 ;
        RECT 104.200 60.800 104.600 63.100 ;
        RECT 105.800 60.800 106.200 63.100 ;
        RECT 108.600 60.800 109.000 65.000 ;
        RECT 110.200 60.800 110.600 63.100 ;
        RECT 111.800 60.800 112.200 65.100 ;
        RECT 115.000 60.800 115.400 65.000 ;
        RECT 117.800 60.800 118.200 63.100 ;
        RECT 119.400 60.800 119.800 63.100 ;
        RECT 122.200 60.800 122.600 65.100 ;
        RECT 123.800 60.800 124.200 65.100 ;
        RECT 125.400 60.800 125.800 65.100 ;
        RECT 127.000 60.800 127.400 65.100 ;
        RECT 128.600 60.800 129.000 65.100 ;
        RECT 130.200 60.800 130.600 65.100 ;
        RECT 131.800 60.800 132.200 65.000 ;
        RECT 134.600 60.800 135.000 63.100 ;
        RECT 136.200 60.800 136.600 63.100 ;
        RECT 139.000 60.800 139.400 65.100 ;
        RECT 140.600 60.800 141.000 65.100 ;
        RECT 142.200 60.800 142.600 65.100 ;
        RECT 143.800 60.800 144.200 65.100 ;
        RECT 145.400 60.800 145.800 65.100 ;
        RECT 147.000 60.800 147.400 65.100 ;
        RECT 150.200 60.800 150.600 64.500 ;
        RECT 152.600 60.800 153.000 64.900 ;
        RECT 154.200 60.800 154.600 63.100 ;
        RECT 155.800 60.800 156.200 64.500 ;
        RECT 158.200 60.800 158.600 64.900 ;
        RECT 159.800 60.800 160.200 63.100 ;
        RECT 160.600 60.800 161.000 63.100 ;
        RECT 162.200 60.800 162.600 63.100 ;
        RECT 163.800 60.800 164.200 62.900 ;
        RECT 165.400 60.800 165.800 63.100 ;
        RECT 166.200 60.800 166.600 65.100 ;
        RECT 167.800 60.800 168.200 63.100 ;
        RECT 169.400 60.800 169.800 63.100 ;
        RECT 170.200 60.800 170.600 65.100 ;
        RECT 173.400 60.800 173.800 65.100 ;
        RECT 174.500 60.800 174.900 63.100 ;
        RECT 176.600 60.800 177.000 65.100 ;
        RECT 179.000 60.800 179.400 65.100 ;
        RECT 180.600 60.800 181.000 65.000 ;
        RECT 183.400 60.800 183.800 63.100 ;
        RECT 185.000 60.800 185.400 63.100 ;
        RECT 187.800 60.800 188.200 65.100 ;
        RECT 190.200 60.800 190.600 64.500 ;
        RECT 192.600 60.800 193.000 64.500 ;
        RECT 0.200 60.200 195.800 60.800 ;
        RECT 0.600 55.900 1.000 60.200 ;
        RECT 2.200 55.900 2.600 60.200 ;
        RECT 3.800 55.900 4.200 60.200 ;
        RECT 5.400 55.900 5.800 60.200 ;
        RECT 7.000 55.900 7.400 60.200 ;
        RECT 7.800 55.900 8.200 60.200 ;
        RECT 11.000 56.100 11.400 60.200 ;
        RECT 13.600 55.900 14.000 60.200 ;
        RECT 15.000 57.900 15.400 60.200 ;
        RECT 16.600 57.900 17.000 60.200 ;
        RECT 17.400 55.900 17.800 60.200 ;
        RECT 19.000 56.500 19.400 60.200 ;
        RECT 20.600 55.900 21.000 60.200 ;
        RECT 23.800 56.100 24.200 60.200 ;
        RECT 26.400 55.900 26.800 60.200 ;
        RECT 27.800 57.900 28.200 60.200 ;
        RECT 29.400 57.900 29.800 60.200 ;
        RECT 31.100 59.900 31.500 60.200 ;
        RECT 31.000 56.600 31.500 59.900 ;
        RECT 34.100 56.600 34.600 60.200 ;
        RECT 35.800 57.900 36.200 60.200 ;
        RECT 37.400 55.900 37.800 60.200 ;
        RECT 39.500 57.900 39.900 60.200 ;
        RECT 40.600 57.900 41.000 60.200 ;
        RECT 42.200 57.900 42.600 60.200 ;
        RECT 43.000 57.900 43.400 60.200 ;
        RECT 46.200 55.900 46.600 60.200 ;
        RECT 48.300 57.900 48.700 60.200 ;
        RECT 49.400 57.900 49.800 60.200 ;
        RECT 51.000 57.900 51.400 60.200 ;
        RECT 52.600 55.900 53.000 60.200 ;
        RECT 55.400 57.900 55.800 60.200 ;
        RECT 57.000 57.900 57.400 60.200 ;
        RECT 59.800 56.000 60.200 60.200 ;
        RECT 62.200 55.900 62.600 60.200 ;
        RECT 65.000 57.900 65.400 60.200 ;
        RECT 66.600 57.900 67.000 60.200 ;
        RECT 69.400 56.000 69.800 60.200 ;
        RECT 71.000 55.900 71.400 60.200 ;
        RECT 73.400 55.900 73.800 60.200 ;
        RECT 76.600 56.100 77.000 60.200 ;
        RECT 79.200 55.900 79.600 60.200 ;
        RECT 81.400 56.500 81.800 60.200 ;
        RECT 86.200 56.500 86.600 60.200 ;
        RECT 87.800 55.900 88.200 60.200 ;
        RECT 90.200 57.900 90.600 60.200 ;
        RECT 91.800 57.900 92.200 60.200 ;
        RECT 92.600 57.900 93.000 60.200 ;
        RECT 96.600 56.900 97.000 60.200 ;
        RECT 103.000 56.500 103.400 60.200 ;
        RECT 107.800 55.900 108.200 60.200 ;
        RECT 108.600 57.900 109.000 60.200 ;
        RECT 110.200 56.100 110.600 60.200 ;
        RECT 114.200 56.500 114.600 60.200 ;
        RECT 116.900 55.900 117.300 60.200 ;
        RECT 119.800 56.500 120.200 60.200 ;
        RECT 123.000 56.500 123.400 60.200 ;
        RECT 125.400 55.900 125.800 60.200 ;
        RECT 128.200 57.900 128.600 60.200 ;
        RECT 129.800 57.900 130.200 60.200 ;
        RECT 132.600 56.000 133.000 60.200 ;
        RECT 135.800 56.500 136.200 60.200 ;
        RECT 139.000 56.500 139.400 60.200 ;
        RECT 140.600 57.900 141.000 60.200 ;
        RECT 142.200 57.900 142.600 60.200 ;
        RECT 143.800 57.900 144.200 60.200 ;
        RECT 145.400 56.500 145.800 60.200 ;
        RECT 149.700 57.900 150.100 60.200 ;
        RECT 151.800 55.900 152.200 60.200 ;
        RECT 152.600 55.900 153.000 60.200 ;
        RECT 155.000 56.600 155.500 60.200 ;
        RECT 158.100 59.900 158.500 60.200 ;
        RECT 158.100 56.600 158.600 59.900 ;
        RECT 161.400 55.900 161.800 60.200 ;
        RECT 163.000 58.100 163.400 60.200 ;
        RECT 164.600 57.900 165.000 60.200 ;
        RECT 165.400 57.900 165.800 60.200 ;
        RECT 167.000 57.900 167.400 60.200 ;
        RECT 167.800 55.900 168.200 60.200 ;
        RECT 170.200 57.900 170.600 60.200 ;
        RECT 171.800 58.100 172.200 60.200 ;
        RECT 173.400 57.900 173.800 60.200 ;
        RECT 175.300 57.900 175.700 60.200 ;
        RECT 177.400 55.900 177.800 60.200 ;
        RECT 178.200 55.900 178.600 60.200 ;
        RECT 180.900 57.900 181.300 60.200 ;
        RECT 183.000 55.900 183.400 60.200 ;
        RECT 184.600 56.000 185.000 60.200 ;
        RECT 187.400 57.900 187.800 60.200 ;
        RECT 189.000 57.900 189.400 60.200 ;
        RECT 191.800 55.900 192.200 60.200 ;
        RECT 194.200 57.900 194.600 60.200 ;
        RECT 1.400 40.800 1.800 44.500 ;
        RECT 3.800 40.800 4.200 45.100 ;
        RECT 6.600 40.800 7.000 43.100 ;
        RECT 8.200 40.800 8.600 43.100 ;
        RECT 11.000 40.800 11.400 45.000 ;
        RECT 14.200 40.800 14.600 45.100 ;
        RECT 15.800 40.800 16.200 45.000 ;
        RECT 18.600 40.800 19.000 43.100 ;
        RECT 20.200 40.800 20.600 43.100 ;
        RECT 23.000 40.800 23.400 45.100 ;
        RECT 25.400 40.800 25.800 45.000 ;
        RECT 28.200 40.800 28.600 43.100 ;
        RECT 29.800 40.800 30.200 43.100 ;
        RECT 32.600 40.800 33.000 45.100 ;
        RECT 39.000 40.800 39.400 44.100 ;
        RECT 41.400 40.800 41.900 44.400 ;
        RECT 44.500 41.100 45.000 44.400 ;
        RECT 44.500 40.800 44.900 41.100 ;
        RECT 48.600 40.800 49.000 45.100 ;
        RECT 51.400 40.800 51.800 43.100 ;
        RECT 53.000 40.800 53.400 43.100 ;
        RECT 55.800 40.800 56.200 45.000 ;
        RECT 57.400 40.800 57.800 45.100 ;
        RECT 59.000 40.800 59.400 45.100 ;
        RECT 60.600 40.800 61.000 45.100 ;
        RECT 62.200 40.800 62.600 45.100 ;
        RECT 63.800 40.800 64.200 45.100 ;
        RECT 65.400 40.800 65.800 44.500 ;
        RECT 67.800 40.800 68.200 43.100 ;
        RECT 69.400 40.800 69.800 45.100 ;
        RECT 72.200 40.800 72.600 43.100 ;
        RECT 73.800 40.800 74.200 43.100 ;
        RECT 76.600 40.800 77.000 45.000 ;
        RECT 78.500 40.800 78.900 43.100 ;
        RECT 80.600 40.800 81.000 45.100 ;
        RECT 81.400 40.800 81.800 43.100 ;
        RECT 83.000 40.800 83.400 43.100 ;
        RECT 85.400 40.800 85.800 45.100 ;
        RECT 87.000 40.800 87.400 45.100 ;
        RECT 87.800 40.800 88.200 45.100 ;
        RECT 90.200 40.800 90.600 43.100 ;
        RECT 91.800 40.800 92.200 43.100 ;
        RECT 92.600 40.800 93.000 45.100 ;
        RECT 100.600 40.800 101.000 44.100 ;
        RECT 103.000 40.800 103.400 43.100 ;
        RECT 104.600 40.800 105.000 44.500 ;
        RECT 107.000 40.800 107.400 44.100 ;
        RECT 113.400 40.800 113.800 44.500 ;
        RECT 117.400 40.800 117.800 44.500 ;
        RECT 120.600 40.800 121.000 45.100 ;
        RECT 123.400 40.800 123.800 43.100 ;
        RECT 125.000 40.800 125.400 43.100 ;
        RECT 127.800 40.800 128.200 45.000 ;
        RECT 130.200 40.800 130.600 45.000 ;
        RECT 133.000 40.800 133.400 43.100 ;
        RECT 134.600 40.800 135.000 43.100 ;
        RECT 137.400 40.800 137.800 45.100 ;
        RECT 139.800 40.800 140.200 45.100 ;
        RECT 142.600 40.800 143.000 43.100 ;
        RECT 144.200 40.800 144.600 43.100 ;
        RECT 147.000 40.800 147.400 45.000 ;
        RECT 150.200 40.800 150.600 45.100 ;
        RECT 152.600 40.800 153.000 45.100 ;
        RECT 155.800 40.800 156.200 42.900 ;
        RECT 157.400 40.800 157.800 43.100 ;
        RECT 159.000 40.800 159.400 45.100 ;
        RECT 161.800 40.800 162.200 43.100 ;
        RECT 163.400 40.800 163.800 43.100 ;
        RECT 166.200 40.800 166.600 45.000 ;
        RECT 167.800 40.800 168.200 43.100 ;
        RECT 169.400 40.800 169.800 43.100 ;
        RECT 170.200 40.800 170.600 45.100 ;
        RECT 173.400 40.800 173.800 45.000 ;
        RECT 176.200 40.800 176.600 43.100 ;
        RECT 177.800 40.800 178.200 43.100 ;
        RECT 180.600 40.800 181.000 45.100 ;
        RECT 183.000 40.800 183.400 45.000 ;
        RECT 185.800 40.800 186.200 43.100 ;
        RECT 187.400 40.800 187.800 43.100 ;
        RECT 190.200 40.800 190.600 45.100 ;
        RECT 192.600 40.800 193.000 44.500 ;
        RECT 0.200 40.200 195.800 40.800 ;
        RECT 1.400 35.900 1.800 40.200 ;
        RECT 4.200 37.900 4.600 40.200 ;
        RECT 5.800 37.900 6.200 40.200 ;
        RECT 8.600 36.000 9.000 40.200 ;
        RECT 11.000 35.900 11.400 40.200 ;
        RECT 13.800 37.900 14.200 40.200 ;
        RECT 15.400 37.900 15.800 40.200 ;
        RECT 18.200 36.000 18.600 40.200 ;
        RECT 20.600 36.000 21.000 40.200 ;
        RECT 23.400 37.900 23.800 40.200 ;
        RECT 25.000 37.900 25.400 40.200 ;
        RECT 27.800 35.900 28.200 40.200 ;
        RECT 30.200 35.900 30.600 40.200 ;
        RECT 33.000 37.900 33.400 40.200 ;
        RECT 34.600 37.900 35.000 40.200 ;
        RECT 37.400 36.000 37.800 40.200 ;
        RECT 39.000 37.900 39.400 40.200 ;
        RECT 40.600 36.100 41.000 40.200 ;
        RECT 42.200 35.900 42.600 40.200 ;
        RECT 45.400 35.900 45.800 40.200 ;
        RECT 48.600 36.100 49.000 40.200 ;
        RECT 50.200 37.900 50.600 40.200 ;
        RECT 52.600 35.900 53.000 40.200 ;
        RECT 54.200 35.900 54.600 40.200 ;
        RECT 57.000 37.900 57.400 40.200 ;
        RECT 58.600 37.900 59.000 40.200 ;
        RECT 61.400 36.000 61.800 40.200 ;
        RECT 64.100 35.900 64.500 40.200 ;
        RECT 66.200 37.900 66.600 40.200 ;
        RECT 67.800 35.900 68.200 40.200 ;
        RECT 70.200 37.900 70.600 40.200 ;
        RECT 71.800 37.900 72.200 40.200 ;
        RECT 73.400 36.100 73.800 40.200 ;
        RECT 75.000 37.900 75.400 40.200 ;
        RECT 75.800 35.900 76.200 40.200 ;
        RECT 78.200 37.900 78.600 40.200 ;
        RECT 80.600 36.000 81.000 40.200 ;
        RECT 83.400 37.900 83.800 40.200 ;
        RECT 85.000 37.900 85.400 40.200 ;
        RECT 87.800 35.900 88.200 40.200 ;
        RECT 90.200 36.000 90.600 40.200 ;
        RECT 93.000 37.900 93.400 40.200 ;
        RECT 94.600 37.900 95.000 40.200 ;
        RECT 97.400 35.900 97.800 40.200 ;
        RECT 101.400 36.100 101.800 40.200 ;
        RECT 103.000 37.900 103.400 40.200 ;
        RECT 104.600 36.900 105.000 40.200 ;
        RECT 111.800 35.900 112.200 40.200 ;
        RECT 113.400 35.900 113.800 40.200 ;
        RECT 116.200 37.900 116.600 40.200 ;
        RECT 117.800 37.900 118.200 40.200 ;
        RECT 120.600 36.000 121.000 40.200 ;
        RECT 122.200 35.900 122.600 40.200 ;
        RECT 125.400 35.900 125.800 40.200 ;
        RECT 128.200 37.900 128.600 40.200 ;
        RECT 129.800 37.900 130.200 40.200 ;
        RECT 132.600 36.000 133.000 40.200 ;
        RECT 135.000 36.500 135.400 40.200 ;
        RECT 137.400 36.500 137.800 40.200 ;
        RECT 139.000 35.900 139.400 40.200 ;
        RECT 140.600 35.900 141.000 40.200 ;
        RECT 142.200 35.900 142.600 40.200 ;
        RECT 143.800 35.900 144.200 40.200 ;
        RECT 145.400 35.900 145.800 40.200 ;
        RECT 148.600 36.000 149.000 40.200 ;
        RECT 151.400 37.900 151.800 40.200 ;
        RECT 153.000 37.900 153.400 40.200 ;
        RECT 155.800 35.900 156.200 40.200 ;
        RECT 158.200 36.000 158.600 40.200 ;
        RECT 161.000 37.900 161.400 40.200 ;
        RECT 162.600 37.900 163.000 40.200 ;
        RECT 165.400 35.900 165.800 40.200 ;
        RECT 168.600 36.500 169.000 40.200 ;
        RECT 171.000 35.900 171.400 40.200 ;
        RECT 173.800 37.900 174.200 40.200 ;
        RECT 175.400 37.900 175.800 40.200 ;
        RECT 178.200 36.000 178.600 40.200 ;
        RECT 180.600 36.000 181.000 40.200 ;
        RECT 183.400 37.900 183.800 40.200 ;
        RECT 185.000 37.900 185.400 40.200 ;
        RECT 187.800 35.900 188.200 40.200 ;
        RECT 190.200 36.500 190.600 40.200 ;
        RECT 192.600 36.500 193.000 40.200 ;
        RECT 135.800 35.100 136.200 35.200 ;
        RECT 136.600 35.100 137.000 35.200 ;
        RECT 135.800 34.800 137.000 35.100 ;
        RECT 135.800 34.400 136.200 34.800 ;
        RECT 136.600 34.400 137.000 34.800 ;
        RECT 189.400 34.400 189.800 35.200 ;
        RECT 191.800 25.800 192.200 26.600 ;
        RECT 1.900 20.800 2.300 25.100 ;
        RECT 5.100 20.800 5.500 25.100 ;
        RECT 7.000 20.800 7.400 23.100 ;
        RECT 9.400 20.800 9.800 25.000 ;
        RECT 12.200 20.800 12.600 23.100 ;
        RECT 13.800 20.800 14.200 23.100 ;
        RECT 16.600 20.800 17.000 25.100 ;
        RECT 19.000 20.800 19.400 25.000 ;
        RECT 21.800 20.800 22.200 23.100 ;
        RECT 23.400 20.800 23.800 23.100 ;
        RECT 26.200 20.800 26.600 25.100 ;
        RECT 28.600 20.800 29.000 25.000 ;
        RECT 31.400 20.800 31.800 23.100 ;
        RECT 33.000 20.800 33.400 23.100 ;
        RECT 35.800 20.800 36.200 25.100 ;
        RECT 39.000 20.800 39.400 25.100 ;
        RECT 40.600 20.800 41.000 25.000 ;
        RECT 43.400 20.800 43.800 23.100 ;
        RECT 45.000 20.800 45.400 23.100 ;
        RECT 47.800 20.800 48.200 25.100 ;
        RECT 51.000 20.800 51.400 23.100 ;
        RECT 52.600 20.800 53.000 24.900 ;
        RECT 55.000 20.800 55.400 25.100 ;
        RECT 57.800 20.800 58.200 23.100 ;
        RECT 59.400 20.800 59.800 23.100 ;
        RECT 62.200 20.800 62.600 25.000 ;
        RECT 64.600 20.800 65.000 24.500 ;
        RECT 67.300 20.800 67.700 25.100 ;
        RECT 69.400 20.800 69.800 25.100 ;
        RECT 71.800 20.800 72.200 23.100 ;
        RECT 73.400 20.800 73.800 23.100 ;
        RECT 75.000 20.800 75.400 22.900 ;
        RECT 76.600 20.800 77.000 25.100 ;
        RECT 79.000 20.800 79.400 25.100 ;
        RECT 81.800 20.800 82.200 23.100 ;
        RECT 83.400 20.800 83.800 23.100 ;
        RECT 86.200 20.800 86.600 25.000 ;
        RECT 88.600 20.800 89.000 25.100 ;
        RECT 91.400 20.800 91.800 23.100 ;
        RECT 93.000 20.800 93.400 23.100 ;
        RECT 95.800 20.800 96.200 25.000 ;
        RECT 99.000 20.800 99.400 23.100 ;
        RECT 100.600 20.800 101.000 24.900 ;
        RECT 103.000 20.800 103.400 25.100 ;
        RECT 105.800 20.800 106.200 23.100 ;
        RECT 107.400 20.800 107.800 23.100 ;
        RECT 110.200 20.800 110.600 25.000 ;
        RECT 112.600 20.800 113.000 25.100 ;
        RECT 115.400 20.800 115.800 23.100 ;
        RECT 117.000 20.800 117.400 23.100 ;
        RECT 119.800 20.800 120.200 25.000 ;
        RECT 121.400 20.800 121.800 23.100 ;
        RECT 123.000 20.800 123.400 25.100 ;
        RECT 124.600 20.800 125.000 25.100 ;
        RECT 126.200 20.800 126.600 25.100 ;
        RECT 127.800 20.800 128.200 25.100 ;
        RECT 129.400 20.800 129.800 25.100 ;
        RECT 130.200 20.800 130.600 23.100 ;
        RECT 131.800 20.800 132.200 25.100 ;
        RECT 135.000 20.800 135.400 25.000 ;
        RECT 137.800 20.800 138.200 23.100 ;
        RECT 139.400 20.800 139.800 23.100 ;
        RECT 142.200 20.800 142.600 25.100 ;
        RECT 146.200 20.800 146.600 25.000 ;
        RECT 149.000 20.800 149.400 23.100 ;
        RECT 150.600 20.800 151.000 23.100 ;
        RECT 153.400 20.800 153.800 25.100 ;
        RECT 155.800 20.800 156.200 25.000 ;
        RECT 158.600 20.800 159.000 23.100 ;
        RECT 160.200 20.800 160.600 23.100 ;
        RECT 163.000 20.800 163.400 25.100 ;
        RECT 164.900 20.800 165.300 23.100 ;
        RECT 167.000 20.800 167.400 25.100 ;
        RECT 168.600 20.800 169.000 25.100 ;
        RECT 171.400 20.800 171.800 23.100 ;
        RECT 173.000 20.800 173.400 23.100 ;
        RECT 175.800 20.800 176.200 25.000 ;
        RECT 177.400 20.800 177.800 25.100 ;
        RECT 180.600 20.800 181.000 25.000 ;
        RECT 183.400 20.800 183.800 23.100 ;
        RECT 185.000 20.800 185.400 23.100 ;
        RECT 187.800 20.800 188.200 25.100 ;
        RECT 190.200 20.800 190.600 24.500 ;
        RECT 192.600 20.800 193.000 24.500 ;
        RECT 0.200 20.200 195.800 20.800 ;
        RECT 1.400 16.500 1.800 20.200 ;
        RECT 3.800 15.900 4.200 20.200 ;
        RECT 6.600 17.900 7.000 20.200 ;
        RECT 8.200 17.900 8.600 20.200 ;
        RECT 11.000 16.000 11.400 20.200 ;
        RECT 14.200 15.900 14.600 20.200 ;
        RECT 15.800 16.000 16.200 20.200 ;
        RECT 18.600 17.900 19.000 20.200 ;
        RECT 20.200 17.900 20.600 20.200 ;
        RECT 23.000 15.900 23.400 20.200 ;
        RECT 26.200 15.900 26.600 20.200 ;
        RECT 27.800 16.500 28.200 20.200 ;
        RECT 30.200 17.900 30.600 20.200 ;
        RECT 31.800 17.900 32.200 20.200 ;
        RECT 32.600 15.900 33.000 20.200 ;
        RECT 35.800 15.900 36.200 20.200 ;
        RECT 38.600 17.900 39.000 20.200 ;
        RECT 40.200 17.900 40.600 20.200 ;
        RECT 43.000 16.000 43.400 20.200 ;
        RECT 46.200 17.900 46.600 20.200 ;
        RECT 47.800 16.100 48.200 20.200 ;
        RECT 50.200 15.900 50.600 20.200 ;
        RECT 53.000 17.900 53.400 20.200 ;
        RECT 54.600 17.900 55.000 20.200 ;
        RECT 57.400 16.000 57.800 20.200 ;
        RECT 59.000 15.900 59.400 20.200 ;
        RECT 60.600 15.900 61.000 20.200 ;
        RECT 62.200 15.900 62.600 20.200 ;
        RECT 63.800 15.900 64.200 20.200 ;
        RECT 65.400 15.900 65.800 20.200 ;
        RECT 67.000 16.000 67.400 20.200 ;
        RECT 69.800 17.900 70.200 20.200 ;
        RECT 71.400 17.900 71.800 20.200 ;
        RECT 74.200 15.900 74.600 20.200 ;
        RECT 76.600 16.100 77.000 20.200 ;
        RECT 78.200 17.900 78.600 20.200 ;
        RECT 79.000 17.900 79.400 20.200 ;
        RECT 80.600 17.900 81.000 20.200 ;
        RECT 83.000 15.900 83.400 20.200 ;
        RECT 83.800 17.900 84.200 20.200 ;
        RECT 86.200 16.500 86.600 20.200 ;
        RECT 88.900 17.900 89.300 20.200 ;
        RECT 91.000 15.900 91.400 20.200 ;
        RECT 93.400 15.900 93.800 20.200 ;
        RECT 95.000 16.500 95.400 20.200 ;
        RECT 99.000 16.900 99.400 20.200 ;
        RECT 104.600 17.900 105.000 20.200 ;
        RECT 106.200 17.900 106.600 20.200 ;
        RECT 107.000 15.900 107.400 20.200 ;
        RECT 109.100 17.900 109.500 20.200 ;
        RECT 110.200 15.900 110.600 20.200 ;
        RECT 114.200 16.500 114.600 20.200 ;
        RECT 116.600 15.900 117.000 20.200 ;
        RECT 119.000 15.900 119.400 20.200 ;
        RECT 120.600 17.900 121.000 20.200 ;
        RECT 122.200 15.900 122.600 20.200 ;
        RECT 125.000 17.900 125.400 20.200 ;
        RECT 126.600 17.900 127.000 20.200 ;
        RECT 129.400 16.000 129.800 20.200 ;
        RECT 131.000 15.900 131.400 20.200 ;
        RECT 133.700 17.900 134.100 20.200 ;
        RECT 135.800 15.900 136.200 20.200 ;
        RECT 136.600 15.900 137.000 20.200 ;
        RECT 138.700 17.900 139.100 20.200 ;
        RECT 140.600 16.500 141.000 20.200 ;
        RECT 143.800 16.000 144.200 20.200 ;
        RECT 146.600 17.900 147.000 20.200 ;
        RECT 148.200 17.900 148.600 20.200 ;
        RECT 151.000 15.900 151.400 20.200 ;
        RECT 154.200 15.900 154.600 20.200 ;
        RECT 156.900 15.900 157.300 20.200 ;
        RECT 159.800 16.000 160.200 20.200 ;
        RECT 162.600 17.900 163.000 20.200 ;
        RECT 164.200 17.900 164.600 20.200 ;
        RECT 167.000 15.900 167.400 20.200 ;
        RECT 168.600 17.900 169.000 20.200 ;
        RECT 170.200 17.900 170.600 20.200 ;
        RECT 172.600 16.500 173.000 20.200 ;
        RECT 175.000 15.900 175.400 20.200 ;
        RECT 175.800 17.900 176.200 20.200 ;
        RECT 177.400 17.900 177.800 20.200 ;
        RECT 178.500 17.900 178.900 20.200 ;
        RECT 180.600 15.900 181.000 20.200 ;
        RECT 183.000 15.900 183.400 20.200 ;
        RECT 183.800 17.900 184.200 20.200 ;
        RECT 186.200 16.000 186.600 20.200 ;
        RECT 189.000 17.900 189.400 20.200 ;
        RECT 190.600 17.900 191.000 20.200 ;
        RECT 193.400 15.900 193.800 20.200 ;
        RECT 0.600 0.800 1.000 3.100 ;
        RECT 2.200 0.800 2.600 5.100 ;
        RECT 4.300 0.800 4.700 3.100 ;
        RECT 7.000 0.800 7.400 5.100 ;
        RECT 12.600 0.800 13.000 4.100 ;
        RECT 15.800 0.800 16.200 5.100 ;
        RECT 16.600 0.800 17.000 3.100 ;
        RECT 18.200 0.800 18.600 3.100 ;
        RECT 19.300 0.800 19.700 3.100 ;
        RECT 21.400 0.800 21.800 5.100 ;
        RECT 22.200 0.800 22.600 5.100 ;
        RECT 23.800 0.800 24.200 5.100 ;
        RECT 31.000 0.800 31.400 4.100 ;
        RECT 32.600 0.800 33.000 3.100 ;
        RECT 34.200 0.800 34.600 3.100 ;
        RECT 35.800 0.800 36.200 5.100 ;
        RECT 38.600 0.800 39.000 3.100 ;
        RECT 40.200 0.800 40.600 3.100 ;
        RECT 43.000 0.800 43.400 5.000 ;
        RECT 46.200 0.800 46.600 5.100 ;
        RECT 48.300 0.800 48.700 3.100 ;
        RECT 49.400 0.800 49.800 5.100 ;
        RECT 51.800 0.800 52.200 3.100 ;
        RECT 53.400 0.800 53.800 5.100 ;
        RECT 55.500 0.800 55.900 3.100 ;
        RECT 57.400 0.800 57.800 4.500 ;
        RECT 59.800 0.800 60.200 4.500 ;
        RECT 62.200 0.800 62.600 3.100 ;
        RECT 63.800 0.800 64.200 3.100 ;
        RECT 65.400 0.800 65.800 5.000 ;
        RECT 68.200 0.800 68.600 3.100 ;
        RECT 69.800 0.800 70.200 3.100 ;
        RECT 72.600 0.800 73.000 5.100 ;
        RECT 74.200 0.800 74.600 3.100 ;
        RECT 76.600 0.800 77.000 4.500 ;
        RECT 80.300 0.800 80.700 5.100 ;
        RECT 82.200 0.800 82.600 3.100 ;
        RECT 83.800 0.800 84.200 3.100 ;
        RECT 85.400 0.800 85.800 2.900 ;
        RECT 87.000 0.800 87.400 3.100 ;
        RECT 88.600 0.800 89.000 3.100 ;
        RECT 90.200 0.800 90.600 5.000 ;
        RECT 93.000 0.800 93.400 3.100 ;
        RECT 94.600 0.800 95.000 3.100 ;
        RECT 97.400 0.800 97.800 5.100 ;
        RECT 100.600 0.800 101.000 5.100 ;
        RECT 103.000 0.800 103.400 3.100 ;
        RECT 104.600 0.800 105.000 3.100 ;
        RECT 106.200 0.800 106.600 4.900 ;
        RECT 107.800 0.800 108.200 3.100 ;
        RECT 109.400 0.800 109.800 5.100 ;
        RECT 112.200 0.800 112.600 3.100 ;
        RECT 113.800 0.800 114.200 3.100 ;
        RECT 116.600 0.800 117.000 5.000 ;
        RECT 118.200 0.800 118.600 3.100 ;
        RECT 119.800 0.800 120.200 3.100 ;
        RECT 122.200 0.800 122.600 5.100 ;
        RECT 123.000 0.800 123.400 5.100 ;
        RECT 125.100 0.800 125.500 3.100 ;
        RECT 126.200 0.800 126.600 3.100 ;
        RECT 127.800 0.800 128.200 3.100 ;
        RECT 129.400 0.800 129.800 5.000 ;
        RECT 132.200 0.800 132.600 3.100 ;
        RECT 133.800 0.800 134.200 3.100 ;
        RECT 136.600 0.800 137.000 5.100 ;
        RECT 138.200 0.800 138.600 3.100 ;
        RECT 139.800 0.800 140.200 4.900 ;
        RECT 142.200 0.800 142.600 5.000 ;
        RECT 145.000 0.800 145.400 3.100 ;
        RECT 146.600 0.800 147.000 3.100 ;
        RECT 149.400 0.800 149.800 5.100 ;
        RECT 153.400 0.800 153.800 5.100 ;
        RECT 156.200 0.800 156.600 3.100 ;
        RECT 157.800 0.800 158.200 3.100 ;
        RECT 160.600 0.800 161.000 5.000 ;
        RECT 162.200 0.800 162.600 5.100 ;
        RECT 165.400 0.800 165.800 4.500 ;
        RECT 167.000 0.800 167.400 5.100 ;
        RECT 169.100 0.800 169.500 3.100 ;
        RECT 170.200 0.800 170.600 5.100 ;
        RECT 173.400 0.800 173.800 5.100 ;
        RECT 176.200 0.800 176.600 3.100 ;
        RECT 177.800 0.800 178.200 3.100 ;
        RECT 180.600 0.800 181.000 5.000 ;
        RECT 183.800 0.800 184.200 5.100 ;
        RECT 185.400 0.800 185.800 5.000 ;
        RECT 188.200 0.800 188.600 3.100 ;
        RECT 189.800 0.800 190.200 3.100 ;
        RECT 192.600 0.800 193.000 5.100 ;
        RECT 0.200 0.200 195.800 0.800 ;
      LAYER via1 ;
        RECT 131.800 163.800 132.200 164.200 ;
        RECT 174.200 163.800 174.600 164.200 ;
        RECT 188.600 163.800 189.000 164.200 ;
        RECT 191.000 163.800 191.400 164.200 ;
        RECT 45.800 160.300 46.200 160.700 ;
        RECT 46.500 160.300 46.900 160.700 ;
        RECT 148.200 160.300 148.600 160.700 ;
        RECT 148.900 160.300 149.300 160.700 ;
        RECT 179.000 156.800 179.400 157.200 ;
        RECT 179.800 154.800 180.200 155.200 ;
        RECT 192.600 154.800 193.000 155.200 ;
        RECT 45.800 140.300 46.200 140.700 ;
        RECT 46.500 140.300 46.900 140.700 ;
        RECT 148.200 140.300 148.600 140.700 ;
        RECT 148.900 140.300 149.300 140.700 ;
        RECT 45.800 120.300 46.200 120.700 ;
        RECT 46.500 120.300 46.900 120.700 ;
        RECT 148.200 120.300 148.600 120.700 ;
        RECT 148.900 120.300 149.300 120.700 ;
        RECT 45.800 100.300 46.200 100.700 ;
        RECT 46.500 100.300 46.900 100.700 ;
        RECT 148.200 100.300 148.600 100.700 ;
        RECT 148.900 100.300 149.300 100.700 ;
        RECT 187.800 83.800 188.200 84.200 ;
        RECT 45.800 80.300 46.200 80.700 ;
        RECT 46.500 80.300 46.900 80.700 ;
        RECT 148.200 80.300 148.600 80.700 ;
        RECT 148.900 80.300 149.300 80.700 ;
        RECT 150.200 74.800 150.600 75.200 ;
        RECT 150.200 63.800 150.600 64.200 ;
        RECT 190.200 63.800 190.600 64.200 ;
        RECT 45.800 60.300 46.200 60.700 ;
        RECT 46.500 60.300 46.900 60.700 ;
        RECT 148.200 60.300 148.600 60.700 ;
        RECT 148.900 60.300 149.300 60.700 ;
        RECT 191.800 59.800 192.200 60.200 ;
        RECT 45.800 40.300 46.200 40.700 ;
        RECT 46.500 40.300 46.900 40.700 ;
        RECT 148.200 40.300 148.600 40.700 ;
        RECT 148.900 40.300 149.300 40.700 ;
        RECT 135.000 36.800 135.400 37.200 ;
        RECT 190.200 36.800 190.600 37.200 ;
        RECT 189.400 34.800 189.800 35.200 ;
        RECT 192.600 23.800 193.000 24.200 ;
        RECT 45.800 20.300 46.200 20.700 ;
        RECT 46.500 20.300 46.900 20.700 ;
        RECT 148.200 20.300 148.600 20.700 ;
        RECT 148.900 20.300 149.300 20.700 ;
        RECT 45.800 0.300 46.200 0.700 ;
        RECT 46.500 0.300 46.900 0.700 ;
        RECT 148.200 0.300 148.600 0.700 ;
        RECT 148.900 0.300 149.300 0.700 ;
      LAYER metal2 ;
        RECT 132.600 165.800 133.000 166.200 ;
        RECT 173.400 165.800 173.800 166.200 ;
        RECT 187.800 165.800 188.200 166.200 ;
        RECT 190.200 165.800 190.600 166.200 ;
        RECT 131.800 164.100 132.200 164.200 ;
        RECT 132.600 164.100 132.900 165.800 ;
        RECT 131.800 163.800 132.900 164.100 ;
        RECT 173.400 164.100 173.700 165.800 ;
        RECT 174.200 164.100 174.600 164.200 ;
        RECT 173.400 163.800 174.600 164.100 ;
        RECT 187.800 164.100 188.100 165.800 ;
        RECT 188.600 164.100 189.000 164.200 ;
        RECT 187.800 163.800 189.000 164.100 ;
        RECT 190.200 164.100 190.500 165.800 ;
        RECT 191.000 164.100 191.400 164.200 ;
        RECT 190.200 163.800 191.400 164.100 ;
        RECT 192.600 160.800 193.000 161.200 ;
        RECT 45.600 160.300 47.200 160.700 ;
        RECT 148.000 160.300 149.600 160.700 ;
        RECT 179.000 157.100 179.400 157.200 ;
        RECT 179.000 156.800 180.100 157.100 ;
        RECT 179.800 155.200 180.100 156.800 ;
        RECT 192.600 155.200 192.900 160.800 ;
        RECT 179.800 154.800 180.200 155.200 ;
        RECT 192.600 155.100 193.000 155.200 ;
        RECT 191.800 154.800 193.000 155.100 ;
        RECT 191.800 146.200 192.100 154.800 ;
        RECT 191.800 145.800 192.200 146.200 ;
        RECT 45.600 140.300 47.200 140.700 ;
        RECT 148.000 140.300 149.600 140.700 ;
        RECT 45.600 120.300 47.200 120.700 ;
        RECT 148.000 120.300 149.600 120.700 ;
        RECT 45.600 100.300 47.200 100.700 ;
        RECT 148.000 100.300 149.600 100.700 ;
        RECT 188.600 85.800 189.000 86.200 ;
        RECT 187.800 84.100 188.200 84.200 ;
        RECT 188.600 84.100 188.900 85.800 ;
        RECT 187.800 83.800 188.900 84.100 ;
        RECT 45.600 80.300 47.200 80.700 ;
        RECT 148.000 80.300 149.600 80.700 ;
        RECT 150.200 74.800 150.600 75.200 ;
        RECT 150.200 64.200 150.500 74.800 ;
        RECT 189.400 65.800 189.800 66.200 ;
        RECT 191.800 65.800 192.200 66.200 ;
        RECT 150.200 63.800 150.600 64.200 ;
        RECT 189.400 64.100 189.700 65.800 ;
        RECT 190.200 64.100 190.600 64.200 ;
        RECT 189.400 63.800 190.600 64.100 ;
        RECT 45.600 60.300 47.200 60.700 ;
        RECT 148.000 60.300 149.600 60.700 ;
        RECT 191.800 60.200 192.100 65.800 ;
        RECT 191.800 59.800 192.200 60.200 ;
        RECT 45.600 40.300 47.200 40.700 ;
        RECT 148.000 40.300 149.600 40.700 ;
        RECT 135.000 37.100 135.400 37.200 ;
        RECT 190.200 37.100 190.600 37.200 ;
        RECT 135.000 36.800 136.100 37.100 ;
        RECT 135.800 35.200 136.100 36.800 ;
        RECT 189.400 36.800 190.600 37.100 ;
        RECT 189.400 35.200 189.700 36.800 ;
        RECT 135.800 34.800 136.200 35.200 ;
        RECT 189.400 34.800 189.800 35.200 ;
        RECT 191.800 25.800 192.200 26.200 ;
        RECT 191.800 24.100 192.100 25.800 ;
        RECT 192.600 24.100 193.000 24.200 ;
        RECT 191.800 23.800 193.000 24.100 ;
        RECT 45.600 20.300 47.200 20.700 ;
        RECT 148.000 20.300 149.600 20.700 ;
        RECT 45.600 0.300 47.200 0.700 ;
        RECT 148.000 0.300 149.600 0.700 ;
      LAYER via2 ;
        RECT 45.800 160.300 46.200 160.700 ;
        RECT 46.500 160.300 46.900 160.700 ;
        RECT 148.200 160.300 148.600 160.700 ;
        RECT 148.900 160.300 149.300 160.700 ;
        RECT 45.800 140.300 46.200 140.700 ;
        RECT 46.500 140.300 46.900 140.700 ;
        RECT 148.200 140.300 148.600 140.700 ;
        RECT 148.900 140.300 149.300 140.700 ;
        RECT 45.800 120.300 46.200 120.700 ;
        RECT 46.500 120.300 46.900 120.700 ;
        RECT 148.200 120.300 148.600 120.700 ;
        RECT 148.900 120.300 149.300 120.700 ;
        RECT 45.800 100.300 46.200 100.700 ;
        RECT 46.500 100.300 46.900 100.700 ;
        RECT 148.200 100.300 148.600 100.700 ;
        RECT 148.900 100.300 149.300 100.700 ;
        RECT 45.800 80.300 46.200 80.700 ;
        RECT 46.500 80.300 46.900 80.700 ;
        RECT 148.200 80.300 148.600 80.700 ;
        RECT 148.900 80.300 149.300 80.700 ;
        RECT 45.800 60.300 46.200 60.700 ;
        RECT 46.500 60.300 46.900 60.700 ;
        RECT 148.200 60.300 148.600 60.700 ;
        RECT 148.900 60.300 149.300 60.700 ;
        RECT 45.800 40.300 46.200 40.700 ;
        RECT 46.500 40.300 46.900 40.700 ;
        RECT 148.200 40.300 148.600 40.700 ;
        RECT 148.900 40.300 149.300 40.700 ;
        RECT 45.800 20.300 46.200 20.700 ;
        RECT 46.500 20.300 46.900 20.700 ;
        RECT 148.200 20.300 148.600 20.700 ;
        RECT 148.900 20.300 149.300 20.700 ;
        RECT 45.800 0.300 46.200 0.700 ;
        RECT 46.500 0.300 46.900 0.700 ;
        RECT 148.200 0.300 148.600 0.700 ;
        RECT 148.900 0.300 149.300 0.700 ;
      LAYER metal3 ;
        RECT 45.600 160.300 47.200 160.700 ;
        RECT 148.000 160.300 149.600 160.700 ;
        RECT 45.600 140.300 47.200 140.700 ;
        RECT 148.000 140.300 149.600 140.700 ;
        RECT 45.600 120.300 47.200 120.700 ;
        RECT 148.000 120.300 149.600 120.700 ;
        RECT 45.600 100.300 47.200 100.700 ;
        RECT 148.000 100.300 149.600 100.700 ;
        RECT 45.600 80.300 47.200 80.700 ;
        RECT 148.000 80.300 149.600 80.700 ;
        RECT 45.600 60.300 47.200 60.700 ;
        RECT 148.000 60.300 149.600 60.700 ;
        RECT 45.600 40.300 47.200 40.700 ;
        RECT 148.000 40.300 149.600 40.700 ;
        RECT 45.600 20.300 47.200 20.700 ;
        RECT 148.000 20.300 149.600 20.700 ;
        RECT 45.600 0.300 47.200 0.700 ;
        RECT 148.000 0.300 149.600 0.700 ;
      LAYER via3 ;
        RECT 45.800 160.300 46.200 160.700 ;
        RECT 46.600 160.300 47.000 160.700 ;
        RECT 148.200 160.300 148.600 160.700 ;
        RECT 149.000 160.300 149.400 160.700 ;
        RECT 45.800 140.300 46.200 140.700 ;
        RECT 46.600 140.300 47.000 140.700 ;
        RECT 148.200 140.300 148.600 140.700 ;
        RECT 149.000 140.300 149.400 140.700 ;
        RECT 45.800 120.300 46.200 120.700 ;
        RECT 46.600 120.300 47.000 120.700 ;
        RECT 148.200 120.300 148.600 120.700 ;
        RECT 149.000 120.300 149.400 120.700 ;
        RECT 45.800 100.300 46.200 100.700 ;
        RECT 46.600 100.300 47.000 100.700 ;
        RECT 148.200 100.300 148.600 100.700 ;
        RECT 149.000 100.300 149.400 100.700 ;
        RECT 45.800 80.300 46.200 80.700 ;
        RECT 46.600 80.300 47.000 80.700 ;
        RECT 148.200 80.300 148.600 80.700 ;
        RECT 149.000 80.300 149.400 80.700 ;
        RECT 45.800 60.300 46.200 60.700 ;
        RECT 46.600 60.300 47.000 60.700 ;
        RECT 148.200 60.300 148.600 60.700 ;
        RECT 149.000 60.300 149.400 60.700 ;
        RECT 45.800 40.300 46.200 40.700 ;
        RECT 46.600 40.300 47.000 40.700 ;
        RECT 148.200 40.300 148.600 40.700 ;
        RECT 149.000 40.300 149.400 40.700 ;
        RECT 45.800 20.300 46.200 20.700 ;
        RECT 46.600 20.300 47.000 20.700 ;
        RECT 148.200 20.300 148.600 20.700 ;
        RECT 149.000 20.300 149.400 20.700 ;
        RECT 45.800 0.300 46.200 0.700 ;
        RECT 46.600 0.300 47.000 0.700 ;
        RECT 148.200 0.300 148.600 0.700 ;
        RECT 149.000 0.300 149.400 0.700 ;
      LAYER metal4 ;
        RECT 45.600 160.300 47.200 160.700 ;
        RECT 148.000 160.300 149.600 160.700 ;
        RECT 45.600 140.300 47.200 140.700 ;
        RECT 148.000 140.300 149.600 140.700 ;
        RECT 45.600 120.300 47.200 120.700 ;
        RECT 148.000 120.300 149.600 120.700 ;
        RECT 45.600 100.300 47.200 100.700 ;
        RECT 148.000 100.300 149.600 100.700 ;
        RECT 45.600 80.300 47.200 80.700 ;
        RECT 148.000 80.300 149.600 80.700 ;
        RECT 45.600 60.300 47.200 60.700 ;
        RECT 148.000 60.300 149.600 60.700 ;
        RECT 45.600 40.300 47.200 40.700 ;
        RECT 148.000 40.300 149.600 40.700 ;
        RECT 45.600 20.300 47.200 20.700 ;
        RECT 148.000 20.300 149.600 20.700 ;
        RECT 45.600 0.300 47.200 0.700 ;
        RECT 148.000 0.300 149.600 0.700 ;
      LAYER via4 ;
        RECT 45.800 160.300 46.200 160.700 ;
        RECT 46.500 160.300 46.900 160.700 ;
        RECT 148.200 160.300 148.600 160.700 ;
        RECT 148.900 160.300 149.300 160.700 ;
        RECT 45.800 140.300 46.200 140.700 ;
        RECT 46.500 140.300 46.900 140.700 ;
        RECT 148.200 140.300 148.600 140.700 ;
        RECT 148.900 140.300 149.300 140.700 ;
        RECT 45.800 120.300 46.200 120.700 ;
        RECT 46.500 120.300 46.900 120.700 ;
        RECT 148.200 120.300 148.600 120.700 ;
        RECT 148.900 120.300 149.300 120.700 ;
        RECT 45.800 100.300 46.200 100.700 ;
        RECT 46.500 100.300 46.900 100.700 ;
        RECT 148.200 100.300 148.600 100.700 ;
        RECT 148.900 100.300 149.300 100.700 ;
        RECT 45.800 80.300 46.200 80.700 ;
        RECT 46.500 80.300 46.900 80.700 ;
        RECT 148.200 80.300 148.600 80.700 ;
        RECT 148.900 80.300 149.300 80.700 ;
        RECT 45.800 60.300 46.200 60.700 ;
        RECT 46.500 60.300 46.900 60.700 ;
        RECT 148.200 60.300 148.600 60.700 ;
        RECT 148.900 60.300 149.300 60.700 ;
        RECT 45.800 40.300 46.200 40.700 ;
        RECT 46.500 40.300 46.900 40.700 ;
        RECT 148.200 40.300 148.600 40.700 ;
        RECT 148.900 40.300 149.300 40.700 ;
        RECT 45.800 20.300 46.200 20.700 ;
        RECT 46.500 20.300 46.900 20.700 ;
        RECT 148.200 20.300 148.600 20.700 ;
        RECT 148.900 20.300 149.300 20.700 ;
        RECT 45.800 0.300 46.200 0.700 ;
        RECT 46.500 0.300 46.900 0.700 ;
        RECT 148.200 0.300 148.600 0.700 ;
        RECT 148.900 0.300 149.300 0.700 ;
      LAYER metal5 ;
        RECT 45.600 160.200 47.200 160.700 ;
        RECT 148.000 160.200 149.600 160.700 ;
        RECT 45.600 140.200 47.200 140.700 ;
        RECT 148.000 140.200 149.600 140.700 ;
        RECT 45.600 120.200 47.200 120.700 ;
        RECT 148.000 120.200 149.600 120.700 ;
        RECT 45.600 100.200 47.200 100.700 ;
        RECT 148.000 100.200 149.600 100.700 ;
        RECT 45.600 80.200 47.200 80.700 ;
        RECT 148.000 80.200 149.600 80.700 ;
        RECT 45.600 60.200 47.200 60.700 ;
        RECT 148.000 60.200 149.600 60.700 ;
        RECT 45.600 40.200 47.200 40.700 ;
        RECT 148.000 40.200 149.600 40.700 ;
        RECT 45.600 20.200 47.200 20.700 ;
        RECT 148.000 20.200 149.600 20.700 ;
        RECT 45.600 0.200 47.200 0.700 ;
        RECT 148.000 0.200 149.600 0.700 ;
      LAYER via5 ;
        RECT 46.600 160.200 47.100 160.700 ;
        RECT 149.000 160.200 149.500 160.700 ;
        RECT 46.600 140.200 47.100 140.700 ;
        RECT 149.000 140.200 149.500 140.700 ;
        RECT 46.600 120.200 47.100 120.700 ;
        RECT 149.000 120.200 149.500 120.700 ;
        RECT 46.600 100.200 47.100 100.700 ;
        RECT 149.000 100.200 149.500 100.700 ;
        RECT 46.600 80.200 47.100 80.700 ;
        RECT 149.000 80.200 149.500 80.700 ;
        RECT 46.600 60.200 47.100 60.700 ;
        RECT 149.000 60.200 149.500 60.700 ;
        RECT 46.600 40.200 47.100 40.700 ;
        RECT 149.000 40.200 149.500 40.700 ;
        RECT 46.600 20.200 47.100 20.700 ;
        RECT 149.000 20.200 149.500 20.700 ;
        RECT 46.600 0.200 47.100 0.700 ;
        RECT 149.000 0.200 149.500 0.700 ;
      LAYER metal6 ;
        RECT 45.600 -3.000 47.200 173.000 ;
        RECT 148.000 -3.000 149.600 173.000 ;
    END
  END vdd
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.200 170.200 195.800 170.800 ;
        RECT 1.400 167.900 1.800 170.200 ;
        RECT 3.800 167.900 4.200 170.200 ;
        RECT 5.400 168.900 5.800 170.200 ;
        RECT 7.000 168.900 7.400 170.200 ;
        RECT 8.600 168.900 9.000 170.200 ;
        RECT 10.200 168.300 10.600 170.200 ;
        RECT 12.600 168.900 13.000 170.200 ;
        RECT 14.700 167.900 15.100 170.200 ;
        RECT 16.600 167.900 17.000 170.200 ;
        RECT 18.200 168.900 18.600 170.200 ;
        RECT 19.800 168.900 20.200 170.200 ;
        RECT 21.400 167.900 21.800 170.200 ;
        RECT 23.800 168.000 24.200 170.200 ;
        RECT 26.600 168.900 27.000 170.200 ;
        RECT 28.200 168.900 28.700 170.200 ;
        RECT 31.000 167.900 31.400 170.200 ;
        RECT 33.400 168.000 33.800 170.200 ;
        RECT 36.200 168.900 36.600 170.200 ;
        RECT 37.800 168.900 38.300 170.200 ;
        RECT 40.600 167.900 41.000 170.200 ;
        RECT 42.200 168.900 42.600 170.200 ;
        RECT 43.800 168.900 44.200 170.200 ;
        RECT 47.000 167.700 47.400 170.200 ;
        RECT 49.600 167.500 50.000 170.200 ;
        RECT 51.800 168.000 52.200 170.200 ;
        RECT 54.600 168.900 55.000 170.200 ;
        RECT 56.200 168.900 56.700 170.200 ;
        RECT 59.000 167.900 59.400 170.200 ;
        RECT 60.600 168.900 61.000 170.200 ;
        RECT 62.200 168.900 62.600 170.200 ;
        RECT 63.800 168.000 64.200 170.200 ;
        RECT 66.600 168.900 67.000 170.200 ;
        RECT 68.200 168.900 68.700 170.200 ;
        RECT 71.000 167.900 71.400 170.200 ;
        RECT 73.400 168.000 73.800 170.200 ;
        RECT 76.200 168.900 76.600 170.200 ;
        RECT 77.800 168.900 78.300 170.200 ;
        RECT 80.600 167.900 81.000 170.200 ;
        RECT 83.000 167.900 83.400 170.200 ;
        RECT 84.600 168.900 85.000 170.200 ;
        RECT 86.200 168.900 86.600 170.200 ;
        RECT 87.800 167.900 88.200 170.200 ;
        RECT 90.200 168.900 90.600 170.200 ;
        RECT 91.800 168.000 92.200 170.200 ;
        RECT 94.600 168.900 95.000 170.200 ;
        RECT 96.200 168.900 96.700 170.200 ;
        RECT 99.000 167.900 99.400 170.200 ;
        RECT 102.200 168.900 102.600 170.200 ;
        RECT 103.800 168.900 104.200 170.200 ;
        RECT 105.400 167.900 105.800 170.200 ;
        RECT 107.800 168.000 108.200 170.200 ;
        RECT 110.600 168.900 111.000 170.200 ;
        RECT 112.200 168.900 112.700 170.200 ;
        RECT 115.000 167.900 115.400 170.200 ;
        RECT 117.400 167.900 117.800 170.200 ;
        RECT 119.800 167.900 120.200 170.200 ;
        RECT 122.200 168.000 122.600 170.200 ;
        RECT 125.000 168.900 125.400 170.200 ;
        RECT 126.600 168.900 127.100 170.200 ;
        RECT 129.400 167.900 129.800 170.200 ;
        RECT 131.800 167.900 132.200 170.200 ;
        RECT 134.200 167.900 134.600 170.200 ;
        RECT 136.600 167.900 137.000 170.200 ;
        RECT 139.300 168.900 139.800 170.200 ;
        RECT 141.000 168.900 141.400 170.200 ;
        RECT 143.800 168.000 144.200 170.200 ;
        RECT 145.400 168.900 145.800 170.200 ;
        RECT 147.000 168.900 147.400 170.200 ;
        RECT 150.200 167.700 150.600 170.200 ;
        RECT 152.800 167.500 153.200 170.200 ;
        RECT 155.000 168.000 155.400 170.200 ;
        RECT 157.800 168.900 158.200 170.200 ;
        RECT 159.400 168.900 159.900 170.200 ;
        RECT 162.200 167.900 162.600 170.200 ;
        RECT 164.600 167.900 165.000 170.200 ;
        RECT 167.300 168.900 167.800 170.200 ;
        RECT 169.000 168.900 169.400 170.200 ;
        RECT 171.800 168.000 172.200 170.200 ;
        RECT 174.200 167.900 174.600 170.200 ;
        RECT 176.600 168.000 177.000 170.200 ;
        RECT 179.400 168.900 179.800 170.200 ;
        RECT 181.000 168.900 181.500 170.200 ;
        RECT 183.800 167.900 184.200 170.200 ;
        RECT 186.200 167.900 186.600 170.200 ;
        RECT 188.600 167.900 189.000 170.200 ;
        RECT 191.000 167.900 191.400 170.200 ;
        RECT 192.600 168.900 193.000 170.200 ;
        RECT 104.600 165.800 105.000 166.600 ;
        RECT 187.000 165.800 187.400 166.600 ;
        RECT 1.400 150.800 1.800 153.000 ;
        RECT 4.200 150.800 4.600 152.100 ;
        RECT 5.800 150.800 6.300 152.100 ;
        RECT 8.600 150.800 9.000 153.100 ;
        RECT 10.800 150.800 11.200 153.500 ;
        RECT 13.400 150.800 13.800 153.300 ;
        RECT 15.600 150.800 16.000 153.500 ;
        RECT 18.200 150.800 18.600 153.300 ;
        RECT 20.400 150.800 20.800 153.500 ;
        RECT 23.000 150.800 23.400 153.300 ;
        RECT 25.200 150.800 25.600 153.500 ;
        RECT 27.800 150.800 28.200 153.300 ;
        RECT 30.200 150.800 30.600 153.000 ;
        RECT 33.000 150.800 33.400 152.100 ;
        RECT 34.600 150.800 35.100 152.100 ;
        RECT 37.400 150.800 37.800 153.100 ;
        RECT 39.800 150.800 40.200 153.100 ;
        RECT 42.500 150.800 43.000 152.100 ;
        RECT 44.200 150.800 44.600 152.100 ;
        RECT 47.000 150.800 47.400 153.000 ;
        RECT 51.000 150.800 51.400 152.100 ;
        RECT 52.600 150.800 53.000 153.000 ;
        RECT 55.400 150.800 55.800 152.100 ;
        RECT 57.000 150.800 57.500 152.100 ;
        RECT 59.800 150.800 60.200 153.100 ;
        RECT 62.200 150.800 62.600 153.000 ;
        RECT 65.000 150.800 65.400 152.100 ;
        RECT 66.600 150.800 67.100 152.100 ;
        RECT 69.400 150.800 69.800 153.100 ;
        RECT 71.800 150.800 72.200 153.000 ;
        RECT 74.600 150.800 75.000 152.100 ;
        RECT 76.200 150.800 76.700 152.100 ;
        RECT 79.000 150.800 79.400 153.100 ;
        RECT 81.400 150.800 81.800 153.000 ;
        RECT 84.200 150.800 84.600 152.100 ;
        RECT 85.800 150.800 86.300 152.100 ;
        RECT 88.600 150.800 89.000 153.100 ;
        RECT 90.800 150.800 91.200 153.500 ;
        RECT 93.400 150.800 93.800 153.300 ;
        RECT 95.300 150.800 95.700 153.100 ;
        RECT 97.400 150.800 97.800 152.100 ;
        RECT 100.600 150.800 101.000 152.700 ;
        RECT 103.000 150.800 103.400 152.100 ;
        RECT 104.600 150.800 105.000 152.100 ;
        RECT 106.200 150.800 106.600 153.100 ;
        RECT 108.600 150.800 109.000 153.100 ;
        RECT 111.000 150.800 111.400 153.300 ;
        RECT 113.600 150.800 114.000 153.500 ;
        RECT 115.800 150.800 116.200 153.100 ;
        RECT 117.400 150.800 117.800 152.100 ;
        RECT 119.000 150.800 119.400 152.100 ;
        RECT 119.800 150.800 120.200 152.100 ;
        RECT 121.900 150.800 122.300 153.100 ;
        RECT 124.600 150.800 125.000 152.700 ;
        RECT 126.200 150.800 126.600 152.100 ;
        RECT 127.800 150.800 128.200 152.100 ;
        RECT 129.400 150.800 129.800 152.100 ;
        RECT 131.000 150.800 131.400 153.100 ;
        RECT 132.600 150.800 133.000 152.100 ;
        RECT 134.200 150.800 134.600 152.100 ;
        RECT 135.800 150.800 136.200 153.000 ;
        RECT 138.600 150.800 139.000 152.100 ;
        RECT 140.200 150.800 140.700 152.100 ;
        RECT 143.000 150.800 143.400 153.100 ;
        RECT 145.200 150.800 145.600 153.500 ;
        RECT 147.800 150.800 148.200 153.300 ;
        RECT 151.000 150.800 151.400 152.100 ;
        RECT 152.600 150.800 153.000 152.100 ;
        RECT 154.200 150.800 154.600 153.100 ;
        RECT 156.900 150.800 157.400 152.100 ;
        RECT 158.600 150.800 159.000 152.100 ;
        RECT 161.400 150.800 161.800 153.000 ;
        RECT 164.100 150.800 164.500 153.000 ;
        RECT 166.200 150.800 166.600 152.100 ;
        RECT 167.800 150.800 168.200 152.100 ;
        RECT 169.200 150.800 169.600 153.500 ;
        RECT 171.800 150.800 172.200 153.300 ;
        RECT 174.200 150.800 174.600 153.300 ;
        RECT 176.800 150.800 177.200 153.500 ;
        RECT 179.000 150.800 179.400 153.100 ;
        RECT 180.600 150.800 181.000 152.100 ;
        RECT 182.200 150.800 182.600 152.100 ;
        RECT 183.800 150.800 184.200 153.100 ;
        RECT 186.500 150.800 187.000 152.100 ;
        RECT 188.200 150.800 188.600 152.100 ;
        RECT 191.000 150.800 191.400 153.000 ;
        RECT 193.400 150.800 193.800 153.100 ;
        RECT 0.200 150.200 195.800 150.800 ;
        RECT 1.400 148.000 1.800 150.200 ;
        RECT 4.200 148.900 4.600 150.200 ;
        RECT 5.800 148.900 6.300 150.200 ;
        RECT 8.600 147.900 9.000 150.200 ;
        RECT 10.200 148.900 10.600 150.200 ;
        RECT 11.800 148.900 12.200 150.200 ;
        RECT 13.400 147.700 13.800 150.200 ;
        RECT 16.000 147.500 16.400 150.200 ;
        RECT 18.200 148.000 18.600 150.200 ;
        RECT 21.000 148.900 21.400 150.200 ;
        RECT 22.600 148.900 23.100 150.200 ;
        RECT 25.400 147.900 25.800 150.200 ;
        RECT 27.800 148.000 28.200 150.200 ;
        RECT 30.600 148.900 31.000 150.200 ;
        RECT 32.200 148.900 32.700 150.200 ;
        RECT 35.000 147.900 35.400 150.200 ;
        RECT 38.200 148.300 38.600 150.200 ;
        RECT 39.800 148.900 40.200 150.200 ;
        RECT 41.900 147.900 42.300 150.200 ;
        RECT 43.000 147.900 43.400 150.200 ;
        RECT 47.000 148.200 47.500 150.200 ;
        RECT 50.100 149.900 50.500 150.200 ;
        RECT 50.100 148.200 50.600 149.900 ;
        RECT 52.100 147.900 52.500 150.200 ;
        RECT 54.200 148.900 54.600 150.200 ;
        RECT 56.600 148.300 57.000 150.200 ;
        RECT 58.200 147.900 58.600 150.200 ;
        RECT 60.100 147.900 60.500 150.200 ;
        RECT 62.200 148.900 62.600 150.200 ;
        RECT 63.800 147.700 64.200 150.200 ;
        RECT 66.400 147.500 66.800 150.200 ;
        RECT 67.800 147.900 68.200 150.200 ;
        RECT 69.400 147.900 69.800 150.200 ;
        RECT 72.600 148.300 73.000 150.200 ;
        RECT 75.000 148.000 75.400 150.200 ;
        RECT 77.800 148.900 78.200 150.200 ;
        RECT 79.400 148.900 79.900 150.200 ;
        RECT 82.200 147.900 82.600 150.200 ;
        RECT 83.800 148.900 84.200 150.200 ;
        RECT 85.400 148.900 85.800 150.200 ;
        RECT 86.500 147.900 86.900 150.200 ;
        RECT 88.600 148.900 89.000 150.200 ;
        RECT 91.000 148.300 91.400 150.200 ;
        RECT 93.200 147.500 93.600 150.200 ;
        RECT 95.800 147.700 96.200 150.200 ;
        RECT 99.800 147.700 100.200 150.200 ;
        RECT 102.400 147.500 102.800 150.200 ;
        RECT 104.600 148.000 105.000 150.200 ;
        RECT 107.400 148.900 107.800 150.200 ;
        RECT 109.000 148.900 109.500 150.200 ;
        RECT 111.800 147.900 112.200 150.200 ;
        RECT 114.200 148.000 114.600 150.200 ;
        RECT 117.000 148.900 117.400 150.200 ;
        RECT 118.600 148.900 119.100 150.200 ;
        RECT 121.400 147.900 121.800 150.200 ;
        RECT 123.000 148.900 123.400 150.200 ;
        RECT 124.600 148.900 125.000 150.200 ;
        RECT 125.400 147.900 125.800 150.200 ;
        RECT 127.000 147.900 127.400 150.200 ;
        RECT 128.600 147.900 129.000 150.200 ;
        RECT 130.200 147.900 130.600 150.200 ;
        RECT 131.800 147.900 132.200 150.200 ;
        RECT 133.400 148.000 133.800 150.200 ;
        RECT 136.200 148.900 136.600 150.200 ;
        RECT 137.800 148.900 138.300 150.200 ;
        RECT 140.600 147.900 141.000 150.200 ;
        RECT 142.200 147.900 142.600 150.200 ;
        RECT 143.800 147.900 144.200 150.200 ;
        RECT 145.400 147.900 145.800 150.200 ;
        RECT 147.000 147.900 147.400 150.200 ;
        RECT 148.600 147.900 149.000 150.200 ;
        RECT 151.800 147.900 152.200 150.200 ;
        RECT 154.500 148.900 155.000 150.200 ;
        RECT 156.200 148.900 156.600 150.200 ;
        RECT 159.000 148.000 159.400 150.200 ;
        RECT 160.600 147.900 161.000 150.200 ;
        RECT 163.800 147.700 164.200 150.200 ;
        RECT 166.400 147.500 166.800 150.200 ;
        RECT 167.800 148.900 168.200 150.200 ;
        RECT 169.400 148.900 169.800 150.200 ;
        RECT 170.200 148.900 170.600 150.200 ;
        RECT 171.800 148.900 172.200 150.200 ;
        RECT 173.400 147.900 173.800 150.200 ;
        RECT 176.100 148.900 176.600 150.200 ;
        RECT 177.800 148.900 178.200 150.200 ;
        RECT 180.600 148.000 181.000 150.200 ;
        RECT 183.000 147.900 183.400 150.200 ;
        RECT 185.700 148.900 186.200 150.200 ;
        RECT 187.400 148.900 187.800 150.200 ;
        RECT 190.200 148.000 190.600 150.200 ;
        RECT 192.600 147.900 193.000 150.200 ;
        RECT 27.000 134.400 27.400 135.200 ;
        RECT 189.400 134.400 189.800 135.200 ;
        RECT 1.400 130.800 1.800 133.000 ;
        RECT 4.200 130.800 4.600 132.100 ;
        RECT 5.800 130.800 6.300 132.100 ;
        RECT 8.600 130.800 9.000 133.100 ;
        RECT 11.000 130.800 11.400 133.100 ;
        RECT 13.700 130.800 14.200 132.100 ;
        RECT 15.400 130.800 15.800 132.100 ;
        RECT 18.200 130.800 18.600 133.000 ;
        RECT 19.800 130.800 20.200 132.100 ;
        RECT 21.400 130.800 21.800 132.100 ;
        RECT 23.000 130.800 23.400 133.300 ;
        RECT 25.600 130.800 26.000 133.500 ;
        RECT 27.800 130.800 28.200 133.100 ;
        RECT 29.400 130.800 29.800 132.100 ;
        RECT 31.000 130.800 31.400 132.100 ;
        RECT 32.400 130.800 32.800 133.500 ;
        RECT 35.000 130.800 35.400 133.300 ;
        RECT 38.200 130.800 38.600 132.700 ;
        RECT 39.800 130.800 40.200 132.100 ;
        RECT 41.900 130.800 42.300 133.100 ;
        RECT 43.000 130.800 43.400 134.100 ;
        RECT 48.600 130.800 49.100 132.800 ;
        RECT 51.700 131.100 52.200 132.800 ;
        RECT 51.700 130.800 52.100 131.100 ;
        RECT 53.400 130.800 53.800 133.100 ;
        RECT 55.000 130.800 55.400 133.100 ;
        RECT 57.400 130.800 57.800 132.700 ;
        RECT 61.400 130.800 61.800 132.700 ;
        RECT 63.000 130.800 63.400 134.100 ;
        RECT 66.200 130.800 66.600 134.100 ;
        RECT 69.400 130.800 69.800 133.100 ;
        RECT 71.800 130.800 72.200 134.100 ;
        RECT 75.800 131.100 76.300 132.800 ;
        RECT 75.900 130.800 76.300 131.100 ;
        RECT 78.900 130.800 79.400 132.800 ;
        RECT 81.400 130.800 81.800 133.300 ;
        RECT 84.000 130.800 84.400 133.500 ;
        RECT 85.700 130.800 86.100 133.100 ;
        RECT 87.800 130.800 88.200 132.100 ;
        RECT 90.200 130.800 90.600 132.700 ;
        RECT 92.400 130.800 92.800 133.500 ;
        RECT 95.000 130.800 95.400 133.300 ;
        RECT 98.200 130.800 98.600 133.100 ;
        RECT 99.800 130.800 100.200 133.100 ;
        RECT 102.200 130.800 102.600 133.300 ;
        RECT 104.800 130.800 105.200 133.500 ;
        RECT 106.800 130.800 107.200 133.500 ;
        RECT 109.400 130.800 109.800 133.300 ;
        RECT 111.000 130.800 111.400 132.100 ;
        RECT 113.200 130.800 113.600 133.500 ;
        RECT 115.800 130.800 116.200 133.300 ;
        RECT 118.200 130.800 118.600 133.300 ;
        RECT 120.800 130.800 121.200 133.500 ;
        RECT 122.800 130.800 123.200 133.500 ;
        RECT 125.400 130.800 125.800 133.300 ;
        RECT 127.800 130.800 128.200 133.300 ;
        RECT 130.400 130.800 130.800 133.500 ;
        RECT 131.800 130.800 132.200 132.100 ;
        RECT 133.900 130.800 134.300 133.100 ;
        RECT 135.800 130.800 136.200 132.700 ;
        RECT 139.000 130.800 139.400 132.900 ;
        RECT 140.600 130.800 141.000 132.100 ;
        RECT 143.000 130.800 143.400 133.100 ;
        RECT 143.800 130.800 144.200 133.100 ;
        RECT 147.800 130.800 148.200 132.700 ;
        RECT 151.000 130.800 151.400 132.100 ;
        RECT 153.400 130.800 153.800 132.700 ;
        RECT 155.800 130.800 156.200 133.100 ;
        RECT 157.700 130.800 158.100 133.100 ;
        RECT 159.800 130.800 160.200 132.100 ;
        RECT 161.400 130.800 161.800 132.700 ;
        RECT 165.400 130.800 165.800 132.700 ;
        RECT 167.000 130.800 167.400 132.100 ;
        RECT 169.100 130.800 169.500 133.100 ;
        RECT 171.000 130.800 171.400 133.100 ;
        RECT 173.700 130.800 174.200 132.100 ;
        RECT 175.400 130.800 175.800 132.100 ;
        RECT 178.200 130.800 178.600 133.000 ;
        RECT 180.600 130.800 181.000 133.000 ;
        RECT 183.400 130.800 183.800 132.100 ;
        RECT 185.000 130.800 185.500 132.100 ;
        RECT 187.800 130.800 188.200 133.100 ;
        RECT 190.200 130.800 190.600 133.100 ;
        RECT 192.600 130.800 193.000 133.100 ;
        RECT 0.200 130.200 195.800 130.800 ;
        RECT 1.400 128.000 1.800 130.200 ;
        RECT 4.200 128.900 4.600 130.200 ;
        RECT 5.800 128.900 6.300 130.200 ;
        RECT 8.600 127.900 9.000 130.200 ;
        RECT 11.000 128.000 11.400 130.200 ;
        RECT 13.800 128.900 14.200 130.200 ;
        RECT 15.400 128.900 15.900 130.200 ;
        RECT 18.200 127.900 18.600 130.200 ;
        RECT 20.600 127.900 21.000 130.200 ;
        RECT 23.300 128.900 23.800 130.200 ;
        RECT 25.000 128.900 25.400 130.200 ;
        RECT 27.800 128.000 28.200 130.200 ;
        RECT 29.400 127.900 29.800 130.200 ;
        RECT 31.000 127.900 31.400 130.200 ;
        RECT 33.400 128.900 33.800 130.200 ;
        RECT 36.600 128.300 37.000 130.200 ;
        RECT 38.200 128.900 38.600 130.200 ;
        RECT 39.800 128.900 40.200 130.200 ;
        RECT 43.000 126.900 43.400 130.200 ;
        RECT 43.800 128.900 44.200 130.200 ;
        RECT 48.600 128.300 49.000 130.200 ;
        RECT 50.200 128.900 50.600 130.200 ;
        RECT 51.800 128.900 52.200 130.200 ;
        RECT 52.600 128.900 53.000 130.200 ;
        RECT 54.200 126.900 54.600 130.200 ;
        RECT 57.400 128.900 57.800 130.200 ;
        RECT 59.000 128.900 59.400 130.200 ;
        RECT 61.400 127.900 61.800 130.200 ;
        RECT 63.800 127.900 64.200 130.200 ;
        RECT 67.000 126.900 67.400 130.200 ;
        RECT 67.800 128.900 68.200 130.200 ;
        RECT 69.400 128.900 69.800 130.200 ;
        RECT 71.000 128.900 71.400 130.200 ;
        RECT 72.600 129.100 73.000 130.200 ;
        RECT 76.600 128.900 77.000 130.200 ;
        RECT 78.200 128.900 78.600 130.200 ;
        RECT 79.800 128.300 80.200 130.200 ;
        RECT 83.800 127.900 84.200 130.200 ;
        RECT 84.600 127.900 85.000 130.200 ;
        RECT 86.200 127.900 86.600 130.200 ;
        RECT 87.000 128.900 87.400 130.200 ;
        RECT 88.600 128.900 89.000 130.200 ;
        RECT 90.200 128.900 90.600 130.200 ;
        RECT 91.800 128.000 92.200 130.200 ;
        RECT 94.600 128.900 95.000 130.200 ;
        RECT 96.200 128.900 96.700 130.200 ;
        RECT 99.000 127.900 99.400 130.200 ;
        RECT 102.200 127.900 102.600 130.200 ;
        RECT 103.800 127.900 104.200 130.200 ;
        RECT 105.400 127.900 105.800 130.200 ;
        RECT 107.000 127.900 107.400 130.200 ;
        RECT 108.600 127.900 109.000 130.200 ;
        RECT 109.400 127.900 109.800 130.200 ;
        RECT 111.000 127.900 111.400 130.200 ;
        RECT 113.400 127.700 113.800 130.200 ;
        RECT 116.000 127.500 116.400 130.200 ;
        RECT 117.400 128.900 117.800 130.200 ;
        RECT 119.000 127.900 119.400 130.200 ;
        RECT 120.600 127.900 121.000 130.200 ;
        RECT 122.200 127.900 122.600 130.200 ;
        RECT 123.800 127.900 124.200 130.200 ;
        RECT 125.400 127.900 125.800 130.200 ;
        RECT 127.000 127.900 127.400 130.200 ;
        RECT 128.600 127.900 129.000 130.200 ;
        RECT 130.200 127.900 130.600 130.200 ;
        RECT 131.800 127.900 132.200 130.200 ;
        RECT 133.400 127.900 133.800 130.200 ;
        RECT 135.000 127.900 135.400 130.200 ;
        RECT 136.600 127.900 137.000 130.200 ;
        RECT 138.200 128.300 138.600 130.200 ;
        RECT 140.600 128.900 141.000 130.200 ;
        RECT 142.700 127.900 143.100 130.200 ;
        RECT 143.800 127.900 144.200 130.200 ;
        RECT 146.200 128.900 146.600 130.200 ;
        RECT 147.800 128.900 148.200 130.200 ;
        RECT 150.200 128.900 150.600 130.200 ;
        RECT 151.800 128.900 152.200 130.200 ;
        RECT 152.900 127.900 153.300 130.200 ;
        RECT 155.000 128.900 155.400 130.200 ;
        RECT 158.200 126.900 158.600 130.200 ;
        RECT 160.600 127.900 161.000 130.200 ;
        RECT 161.400 128.900 161.800 130.200 ;
        RECT 163.000 128.900 163.400 130.200 ;
        RECT 165.400 128.300 165.800 130.200 ;
        RECT 167.800 128.200 168.300 130.200 ;
        RECT 170.900 129.900 171.300 130.200 ;
        RECT 170.900 128.200 171.400 129.900 ;
        RECT 173.400 128.000 173.800 130.200 ;
        RECT 176.200 128.900 176.600 130.200 ;
        RECT 177.800 128.900 178.300 130.200 ;
        RECT 180.600 127.900 181.000 130.200 ;
        RECT 182.800 127.500 183.200 130.200 ;
        RECT 185.400 127.700 185.800 130.200 ;
        RECT 187.000 128.900 187.400 130.200 ;
        RECT 188.600 128.900 189.000 130.200 ;
        RECT 190.200 128.900 190.600 130.200 ;
        RECT 191.800 127.900 192.200 130.200 ;
        RECT 193.400 128.900 193.800 130.200 ;
        RECT 195.000 128.900 195.400 130.200 ;
        RECT 191.800 114.400 192.200 115.200 ;
        RECT 1.400 110.800 1.800 113.000 ;
        RECT 4.200 110.800 4.600 112.100 ;
        RECT 5.800 110.800 6.300 112.100 ;
        RECT 8.600 110.800 9.000 113.100 ;
        RECT 10.200 110.800 10.600 112.100 ;
        RECT 11.800 110.800 12.200 112.100 ;
        RECT 13.900 110.800 14.300 113.000 ;
        RECT 16.600 110.800 17.000 113.100 ;
        RECT 19.300 110.800 19.800 112.100 ;
        RECT 21.000 110.800 21.400 112.100 ;
        RECT 23.800 110.800 24.200 113.000 ;
        RECT 26.200 110.800 26.600 113.000 ;
        RECT 29.000 110.800 29.400 112.100 ;
        RECT 30.600 110.800 31.100 112.100 ;
        RECT 33.400 110.800 33.800 113.100 ;
        RECT 35.800 110.800 36.200 112.700 ;
        RECT 38.200 110.800 38.600 112.100 ;
        RECT 40.300 110.800 40.700 113.100 ;
        RECT 41.400 110.800 41.800 112.100 ;
        RECT 43.000 110.800 43.400 112.100 ;
        RECT 46.200 110.800 46.600 114.100 ;
        RECT 51.000 110.800 51.400 114.100 ;
        RECT 54.200 110.800 54.600 114.100 ;
        RECT 55.800 110.800 56.200 112.100 ;
        RECT 58.200 110.800 58.600 113.100 ;
        RECT 60.600 110.800 61.000 112.700 ;
        RECT 63.000 110.800 63.400 112.100 ;
        RECT 64.900 110.800 65.300 113.000 ;
        RECT 67.000 110.800 67.400 112.100 ;
        RECT 68.600 110.800 69.000 112.100 ;
        RECT 70.200 110.800 70.600 113.000 ;
        RECT 73.000 110.800 73.400 112.100 ;
        RECT 74.600 110.800 75.100 112.100 ;
        RECT 77.400 110.800 77.800 113.100 ;
        RECT 79.800 110.800 80.200 112.100 ;
        RECT 81.400 110.800 81.800 112.700 ;
        RECT 85.400 110.800 85.800 113.100 ;
        RECT 87.000 110.800 87.400 113.300 ;
        RECT 89.600 110.800 90.000 113.500 ;
        RECT 91.000 110.800 91.400 112.100 ;
        RECT 92.600 110.800 93.000 112.100 ;
        RECT 95.800 110.800 96.200 113.000 ;
        RECT 98.600 110.800 99.000 112.100 ;
        RECT 100.200 110.800 100.700 112.100 ;
        RECT 103.000 110.800 103.400 113.100 ;
        RECT 105.400 110.800 105.800 113.100 ;
        RECT 108.100 110.800 108.600 112.100 ;
        RECT 109.800 110.800 110.200 112.100 ;
        RECT 112.600 110.800 113.000 113.000 ;
        RECT 115.000 110.800 115.400 113.000 ;
        RECT 117.800 110.800 118.200 112.100 ;
        RECT 119.400 110.800 119.900 112.100 ;
        RECT 122.200 110.800 122.600 113.100 ;
        RECT 123.800 110.800 124.200 112.100 ;
        RECT 125.400 110.800 125.800 112.100 ;
        RECT 126.800 110.800 127.200 113.500 ;
        RECT 129.400 110.800 129.800 113.300 ;
        RECT 132.600 110.800 133.000 113.100 ;
        RECT 133.400 110.800 133.800 112.100 ;
        RECT 135.000 110.800 135.400 112.100 ;
        RECT 135.800 110.800 136.200 113.100 ;
        RECT 139.800 110.800 140.200 112.700 ;
        RECT 142.200 110.800 142.600 112.100 ;
        RECT 143.800 110.800 144.200 112.100 ;
        RECT 147.000 110.800 147.400 113.000 ;
        RECT 149.800 110.800 150.200 112.100 ;
        RECT 151.400 110.800 151.900 112.100 ;
        RECT 154.200 110.800 154.600 113.100 ;
        RECT 157.100 110.800 157.500 113.000 ;
        RECT 159.800 110.800 160.200 113.000 ;
        RECT 162.600 110.800 163.000 112.100 ;
        RECT 164.200 110.800 164.700 112.100 ;
        RECT 167.000 110.800 167.400 113.100 ;
        RECT 169.400 110.800 169.800 113.000 ;
        RECT 172.200 110.800 172.600 112.100 ;
        RECT 173.800 110.800 174.300 112.100 ;
        RECT 176.600 110.800 177.000 113.100 ;
        RECT 178.800 110.800 179.200 113.500 ;
        RECT 181.400 110.800 181.800 113.300 ;
        RECT 184.600 110.800 185.000 112.700 ;
        RECT 187.000 110.800 187.400 113.100 ;
        RECT 188.900 110.800 189.300 113.100 ;
        RECT 191.000 110.800 191.400 112.100 ;
        RECT 192.600 110.800 193.000 113.100 ;
        RECT 0.200 110.200 195.800 110.800 ;
        RECT 0.600 107.900 1.000 110.200 ;
        RECT 4.600 108.300 5.000 110.200 ;
        RECT 7.000 108.900 7.400 110.200 ;
        RECT 9.100 108.000 9.500 110.200 ;
        RECT 11.000 108.900 11.400 110.200 ;
        RECT 12.600 108.900 13.000 110.200 ;
        RECT 15.800 108.300 16.200 110.200 ;
        RECT 17.400 107.900 17.800 110.200 ;
        RECT 21.400 108.300 21.800 110.200 ;
        RECT 23.800 108.900 24.200 110.200 ;
        RECT 25.500 109.900 25.900 110.200 ;
        RECT 25.400 108.200 25.900 109.900 ;
        RECT 28.500 108.200 29.000 110.200 ;
        RECT 30.200 107.900 30.600 110.200 ;
        RECT 34.200 108.300 34.600 110.200 ;
        RECT 36.600 108.900 37.000 110.200 ;
        RECT 37.400 107.900 37.800 110.200 ;
        RECT 39.800 106.900 40.200 110.200 ;
        RECT 45.400 108.900 45.800 110.200 ;
        RECT 47.000 109.100 47.400 110.200 ;
        RECT 51.000 107.900 51.400 110.200 ;
        RECT 52.600 107.900 53.000 110.200 ;
        RECT 55.000 107.700 55.400 110.200 ;
        RECT 57.600 107.500 58.000 110.200 ;
        RECT 59.000 107.900 59.400 110.200 ;
        RECT 62.200 108.300 62.600 110.200 ;
        RECT 65.400 108.900 65.800 110.200 ;
        RECT 67.000 108.900 67.400 110.200 ;
        RECT 69.100 108.000 69.500 110.200 ;
        RECT 72.600 108.300 73.000 110.200 ;
        RECT 75.000 108.900 75.400 110.200 ;
        RECT 75.800 107.900 76.200 110.200 ;
        RECT 77.400 107.900 77.800 110.200 ;
        RECT 79.000 107.900 79.400 110.200 ;
        RECT 80.600 107.900 81.000 110.200 ;
        RECT 82.200 107.900 82.600 110.200 ;
        RECT 83.800 108.000 84.200 110.200 ;
        RECT 86.600 108.900 87.000 110.200 ;
        RECT 88.200 108.900 88.700 110.200 ;
        RECT 91.000 107.900 91.400 110.200 ;
        RECT 95.000 108.000 95.400 110.200 ;
        RECT 97.800 108.900 98.200 110.200 ;
        RECT 99.400 108.900 99.900 110.200 ;
        RECT 102.200 107.900 102.600 110.200 ;
        RECT 104.600 108.000 105.000 110.200 ;
        RECT 107.400 108.900 107.800 110.200 ;
        RECT 109.000 108.900 109.500 110.200 ;
        RECT 111.800 107.900 112.200 110.200 ;
        RECT 113.400 108.900 113.800 110.200 ;
        RECT 115.000 108.900 115.400 110.200 ;
        RECT 115.800 107.900 116.200 110.200 ;
        RECT 117.400 107.900 117.800 110.200 ;
        RECT 119.000 107.900 119.400 110.200 ;
        RECT 120.600 107.900 121.000 110.200 ;
        RECT 122.200 107.900 122.600 110.200 ;
        RECT 123.800 107.700 124.200 110.200 ;
        RECT 126.400 107.500 126.800 110.200 ;
        RECT 128.600 107.900 129.000 110.200 ;
        RECT 131.300 108.900 131.800 110.200 ;
        RECT 133.000 108.900 133.400 110.200 ;
        RECT 135.800 108.000 136.200 110.200 ;
        RECT 138.200 107.900 138.600 110.200 ;
        RECT 140.900 108.900 141.400 110.200 ;
        RECT 142.600 108.900 143.000 110.200 ;
        RECT 145.400 108.000 145.800 110.200 ;
        RECT 147.000 107.900 147.400 110.200 ;
        RECT 152.600 108.300 153.000 110.200 ;
        RECT 155.000 108.900 155.400 110.200 ;
        RECT 155.800 108.900 156.200 110.200 ;
        RECT 157.400 108.900 157.800 110.200 ;
        RECT 160.600 108.300 161.000 110.200 ;
        RECT 162.200 108.900 162.600 110.200 ;
        RECT 163.800 108.900 164.200 110.200 ;
        RECT 165.700 108.000 166.100 110.200 ;
        RECT 168.600 107.700 169.000 110.200 ;
        RECT 171.200 107.500 171.600 110.200 ;
        RECT 172.600 108.900 173.000 110.200 ;
        RECT 174.200 108.900 174.600 110.200 ;
        RECT 175.000 107.900 175.400 110.200 ;
        RECT 176.600 107.900 177.000 110.200 ;
        RECT 178.200 107.900 178.600 110.200 ;
        RECT 179.800 107.900 180.200 110.200 ;
        RECT 181.400 107.900 181.800 110.200 ;
        RECT 182.800 107.500 183.200 110.200 ;
        RECT 185.400 107.700 185.800 110.200 ;
        RECT 187.800 107.700 188.200 110.200 ;
        RECT 190.400 107.500 190.800 110.200 ;
        RECT 191.800 108.900 192.200 110.200 ;
        RECT 193.400 108.100 193.800 110.200 ;
        RECT 192.600 94.400 193.000 95.200 ;
        RECT 1.400 90.800 1.800 93.100 ;
        RECT 4.600 90.800 5.000 92.700 ;
        RECT 7.000 90.800 7.400 92.100 ;
        RECT 8.600 91.100 9.100 92.800 ;
        RECT 8.700 90.800 9.100 91.100 ;
        RECT 11.700 90.800 12.200 92.800 ;
        RECT 14.200 90.800 14.600 93.000 ;
        RECT 17.000 90.800 17.400 92.100 ;
        RECT 18.600 90.800 19.100 92.100 ;
        RECT 21.400 90.800 21.800 93.100 ;
        RECT 26.200 90.800 26.600 91.900 ;
        RECT 27.800 90.800 28.200 92.100 ;
        RECT 29.400 90.800 29.800 92.100 ;
        RECT 31.500 90.800 31.900 93.100 ;
        RECT 33.400 90.800 33.800 92.700 ;
        RECT 36.600 90.800 37.000 92.700 ;
        RECT 39.000 90.800 39.400 92.100 ;
        RECT 40.600 90.800 41.000 92.100 ;
        RECT 43.000 90.800 43.400 93.100 ;
        RECT 43.800 90.800 44.200 92.100 ;
        RECT 45.900 90.800 46.300 93.100 ;
        RECT 49.400 90.800 49.900 92.800 ;
        RECT 52.500 91.100 53.000 92.800 ;
        RECT 52.500 90.800 52.900 91.100 ;
        RECT 55.800 90.800 56.200 93.100 ;
        RECT 57.400 90.800 57.800 92.100 ;
        RECT 59.000 90.800 59.400 91.900 ;
        RECT 63.800 90.800 64.300 92.800 ;
        RECT 66.900 91.100 67.400 92.800 ;
        RECT 66.900 90.800 67.300 91.100 ;
        RECT 68.600 90.800 69.000 92.100 ;
        RECT 71.000 90.800 71.400 92.700 ;
        RECT 74.200 90.800 74.600 93.300 ;
        RECT 76.800 90.800 77.200 93.500 ;
        RECT 78.200 90.800 78.600 92.100 ;
        RECT 79.800 90.800 80.200 92.100 ;
        RECT 81.400 90.800 81.800 93.300 ;
        RECT 84.000 90.800 84.400 93.500 ;
        RECT 85.400 90.800 85.800 92.100 ;
        RECT 87.000 90.800 87.400 92.100 ;
        RECT 88.600 90.800 89.000 93.000 ;
        RECT 91.400 90.800 91.800 92.100 ;
        RECT 93.000 90.800 93.500 92.100 ;
        RECT 95.800 90.800 96.200 93.100 ;
        RECT 99.000 90.800 99.400 93.100 ;
        RECT 100.600 90.800 101.000 93.100 ;
        RECT 102.200 90.800 102.600 93.100 ;
        RECT 103.800 90.800 104.200 93.100 ;
        RECT 105.400 90.800 105.800 93.100 ;
        RECT 106.200 90.800 106.600 92.100 ;
        RECT 107.800 90.800 108.200 92.100 ;
        RECT 109.400 90.800 109.800 93.300 ;
        RECT 112.000 90.800 112.400 93.500 ;
        RECT 115.000 90.800 115.400 92.700 ;
        RECT 118.200 90.800 118.600 93.100 ;
        RECT 119.800 90.800 120.200 92.100 ;
        RECT 122.200 90.800 122.600 92.700 ;
        RECT 124.600 90.800 125.000 92.100 ;
        RECT 126.200 90.800 126.700 92.800 ;
        RECT 129.300 91.100 129.800 92.800 ;
        RECT 129.300 90.800 129.700 91.100 ;
        RECT 131.800 90.800 132.200 92.100 ;
        RECT 133.400 90.800 133.800 91.900 ;
        RECT 138.200 91.100 138.700 92.800 ;
        RECT 138.300 90.800 138.700 91.100 ;
        RECT 141.300 90.800 141.800 92.800 ;
        RECT 143.800 90.800 144.200 93.000 ;
        RECT 146.600 90.800 147.000 92.100 ;
        RECT 148.200 90.800 148.700 92.100 ;
        RECT 151.000 90.800 151.400 93.100 ;
        RECT 155.000 90.800 155.400 93.000 ;
        RECT 157.800 90.800 158.200 92.100 ;
        RECT 159.400 90.800 159.900 92.100 ;
        RECT 162.200 90.800 162.600 93.100 ;
        RECT 164.600 90.800 165.000 93.100 ;
        RECT 167.300 90.800 167.800 92.100 ;
        RECT 169.000 90.800 169.400 92.100 ;
        RECT 171.800 90.800 172.200 93.000 ;
        RECT 174.200 90.800 174.600 93.000 ;
        RECT 177.000 90.800 177.400 92.100 ;
        RECT 178.600 90.800 179.100 92.100 ;
        RECT 181.400 90.800 181.800 93.100 ;
        RECT 183.800 90.800 184.200 93.100 ;
        RECT 186.500 90.800 187.000 92.100 ;
        RECT 188.200 90.800 188.600 92.100 ;
        RECT 191.000 90.800 191.400 93.000 ;
        RECT 193.400 90.800 193.800 93.100 ;
        RECT 0.200 90.200 195.800 90.800 ;
        RECT 0.600 87.900 1.000 90.200 ;
        RECT 3.600 87.500 4.000 90.200 ;
        RECT 6.200 87.700 6.600 90.200 ;
        RECT 8.600 87.700 9.000 90.200 ;
        RECT 11.200 87.500 11.600 90.200 ;
        RECT 13.400 88.000 13.800 90.200 ;
        RECT 16.200 88.900 16.600 90.200 ;
        RECT 17.800 88.900 18.300 90.200 ;
        RECT 20.600 87.900 21.000 90.200 ;
        RECT 22.200 87.900 22.600 90.200 ;
        RECT 23.800 87.900 24.200 90.200 ;
        RECT 26.200 87.900 26.600 90.200 ;
        RECT 27.800 87.900 28.200 90.200 ;
        RECT 28.600 87.900 29.000 90.200 ;
        RECT 30.200 88.900 30.600 90.200 ;
        RECT 31.800 88.900 32.200 90.200 ;
        RECT 32.600 87.900 33.000 90.200 ;
        RECT 35.000 88.900 35.400 90.200 ;
        RECT 36.600 87.900 37.000 90.200 ;
        RECT 39.000 87.900 39.400 90.200 ;
        RECT 43.000 88.300 43.400 90.200 ;
        RECT 44.600 88.900 45.000 90.200 ;
        RECT 46.200 88.900 46.600 90.200 ;
        RECT 49.500 89.900 49.900 90.200 ;
        RECT 49.400 88.200 49.900 89.900 ;
        RECT 52.500 88.200 53.000 90.200 ;
        RECT 55.800 88.300 56.200 90.200 ;
        RECT 58.200 88.900 58.600 90.200 ;
        RECT 59.000 86.900 59.400 90.200 ;
        RECT 63.000 88.000 63.400 90.200 ;
        RECT 65.800 88.900 66.200 90.200 ;
        RECT 67.400 88.900 67.900 90.200 ;
        RECT 70.200 87.900 70.600 90.200 ;
        RECT 73.400 87.900 73.800 90.200 ;
        RECT 75.000 88.000 75.400 90.200 ;
        RECT 77.800 88.900 78.200 90.200 ;
        RECT 79.400 88.900 79.900 90.200 ;
        RECT 82.200 87.900 82.600 90.200 ;
        RECT 83.800 87.900 84.200 90.200 ;
        RECT 85.400 87.900 85.800 90.200 ;
        RECT 87.800 88.000 88.200 90.200 ;
        RECT 90.600 88.900 91.000 90.200 ;
        RECT 92.200 88.900 92.700 90.200 ;
        RECT 95.000 87.900 95.400 90.200 ;
        RECT 99.000 88.000 99.400 90.200 ;
        RECT 101.800 88.900 102.200 90.200 ;
        RECT 103.400 88.900 103.900 90.200 ;
        RECT 106.200 87.900 106.600 90.200 ;
        RECT 108.600 88.000 109.000 90.200 ;
        RECT 111.400 88.900 111.800 90.200 ;
        RECT 113.000 88.900 113.500 90.200 ;
        RECT 115.800 87.900 116.200 90.200 ;
        RECT 117.400 88.900 117.800 90.200 ;
        RECT 119.000 88.900 119.400 90.200 ;
        RECT 121.400 87.900 121.800 90.200 ;
        RECT 123.000 87.700 123.400 90.200 ;
        RECT 125.600 87.500 126.000 90.200 ;
        RECT 127.800 88.000 128.200 90.200 ;
        RECT 130.600 88.900 131.000 90.200 ;
        RECT 132.200 88.900 132.700 90.200 ;
        RECT 135.000 87.900 135.400 90.200 ;
        RECT 136.600 88.900 137.000 90.200 ;
        RECT 138.200 88.900 138.600 90.200 ;
        RECT 139.600 87.500 140.000 90.200 ;
        RECT 142.200 87.700 142.600 90.200 ;
        RECT 146.200 88.000 146.600 90.200 ;
        RECT 149.000 88.900 149.400 90.200 ;
        RECT 150.600 88.900 151.100 90.200 ;
        RECT 153.400 87.900 153.800 90.200 ;
        RECT 155.800 87.900 156.200 90.200 ;
        RECT 158.200 88.300 158.600 90.200 ;
        RECT 162.200 87.900 162.600 90.200 ;
        RECT 165.400 86.900 165.800 90.200 ;
        RECT 166.200 86.900 166.600 90.200 ;
        RECT 169.400 88.900 169.800 90.200 ;
        RECT 171.000 88.900 171.400 90.200 ;
        RECT 171.800 87.900 172.200 90.200 ;
        RECT 174.200 88.300 174.600 90.200 ;
        RECT 176.600 88.900 177.000 90.200 ;
        RECT 178.200 88.900 178.600 90.200 ;
        RECT 179.000 88.900 179.400 90.200 ;
        RECT 180.600 88.900 181.000 90.200 ;
        RECT 182.200 88.200 182.700 90.200 ;
        RECT 185.300 89.900 185.700 90.200 ;
        RECT 185.300 88.200 185.800 89.900 ;
        RECT 187.800 87.900 188.200 90.200 ;
        RECT 190.200 87.900 190.600 90.200 ;
        RECT 192.600 87.900 193.000 90.200 ;
        RECT 155.000 85.800 155.400 86.600 ;
        RECT 189.400 85.800 189.800 86.600 ;
        RECT 0.600 70.800 1.000 73.100 ;
        RECT 2.200 70.800 2.600 73.100 ;
        RECT 3.800 70.800 4.200 73.100 ;
        RECT 5.400 70.800 5.800 73.100 ;
        RECT 7.000 70.800 7.400 73.100 ;
        RECT 7.800 70.800 8.200 72.100 ;
        RECT 9.400 70.800 9.800 72.100 ;
        RECT 11.000 70.800 11.400 73.000 ;
        RECT 13.800 70.800 14.200 72.100 ;
        RECT 15.400 70.800 15.900 72.100 ;
        RECT 18.200 70.800 18.600 73.100 ;
        RECT 20.600 70.800 21.000 73.100 ;
        RECT 23.300 70.800 23.800 72.100 ;
        RECT 25.000 70.800 25.400 72.100 ;
        RECT 27.800 70.800 28.200 73.000 ;
        RECT 29.400 70.800 29.800 72.100 ;
        RECT 31.000 70.800 31.400 72.100 ;
        RECT 32.600 70.800 33.000 73.000 ;
        RECT 35.400 70.800 35.800 72.100 ;
        RECT 37.000 70.800 37.500 72.100 ;
        RECT 39.800 70.800 40.200 73.100 ;
        RECT 41.400 70.800 41.800 72.100 ;
        RECT 43.000 70.800 43.400 72.100 ;
        RECT 43.800 70.800 44.200 73.100 ;
        RECT 47.800 70.800 48.200 72.100 ;
        RECT 49.400 70.800 49.800 72.100 ;
        RECT 51.000 70.800 51.400 72.100 ;
        RECT 53.400 70.800 53.800 73.100 ;
        RECT 55.800 70.800 56.200 72.700 ;
        RECT 57.400 70.800 57.800 72.100 ;
        RECT 59.000 70.800 59.400 72.900 ;
        RECT 60.900 70.800 61.300 73.100 ;
        RECT 63.000 70.800 63.400 72.100 ;
        RECT 66.200 70.800 66.600 74.100 ;
        RECT 67.800 70.800 68.200 73.000 ;
        RECT 70.600 70.800 71.000 72.100 ;
        RECT 72.200 70.800 72.700 72.100 ;
        RECT 75.000 70.800 75.400 73.100 ;
        RECT 76.900 70.800 77.300 73.100 ;
        RECT 79.000 70.800 79.400 72.100 ;
        RECT 80.600 70.800 81.000 72.700 ;
        RECT 84.600 70.800 85.000 72.700 ;
        RECT 87.800 70.800 88.200 72.700 ;
        RECT 89.400 70.800 89.800 73.100 ;
        RECT 91.000 70.800 91.400 73.100 ;
        RECT 93.200 70.800 93.600 73.500 ;
        RECT 95.800 70.800 96.200 73.300 ;
        RECT 99.800 70.800 100.200 73.100 ;
        RECT 101.400 70.800 101.800 73.100 ;
        RECT 102.200 70.800 102.600 73.100 ;
        RECT 103.800 70.800 104.200 73.100 ;
        RECT 105.400 70.800 105.800 73.100 ;
        RECT 107.000 70.800 107.400 73.100 ;
        RECT 109.700 70.800 110.200 72.100 ;
        RECT 111.400 70.800 111.800 72.100 ;
        RECT 114.200 70.800 114.600 73.000 ;
        RECT 116.600 70.800 117.000 73.100 ;
        RECT 119.300 70.800 119.800 72.100 ;
        RECT 121.000 70.800 121.400 72.100 ;
        RECT 123.800 70.800 124.200 73.000 ;
        RECT 125.400 70.800 125.800 72.100 ;
        RECT 127.000 70.800 127.400 72.100 ;
        RECT 127.800 70.800 128.200 73.100 ;
        RECT 129.400 70.800 129.800 73.100 ;
        RECT 131.000 70.800 131.400 73.100 ;
        RECT 132.600 70.800 133.000 73.100 ;
        RECT 134.200 70.800 134.600 73.100 ;
        RECT 135.000 70.800 135.400 73.100 ;
        RECT 136.600 70.800 137.000 73.100 ;
        RECT 138.200 70.800 138.600 73.100 ;
        RECT 139.800 70.800 140.200 73.100 ;
        RECT 142.500 70.800 143.000 72.100 ;
        RECT 144.200 70.800 144.600 72.100 ;
        RECT 147.000 70.800 147.400 73.000 ;
        RECT 151.000 70.800 151.400 73.100 ;
        RECT 152.600 70.800 153.000 72.100 ;
        RECT 155.000 70.800 155.400 73.100 ;
        RECT 157.700 70.800 158.200 72.100 ;
        RECT 159.400 70.800 159.800 72.100 ;
        RECT 162.200 70.800 162.600 73.000 ;
        RECT 163.800 70.800 164.200 72.100 ;
        RECT 165.400 70.800 165.800 72.100 ;
        RECT 166.200 70.800 166.600 73.100 ;
        RECT 168.600 70.800 169.000 72.100 ;
        RECT 171.800 70.800 172.200 72.700 ;
        RECT 173.400 70.800 173.800 72.100 ;
        RECT 175.000 70.800 175.400 72.100 ;
        RECT 176.600 70.800 177.000 72.100 ;
        RECT 177.400 70.800 177.800 72.100 ;
        RECT 179.500 70.800 179.900 73.100 ;
        RECT 182.200 70.800 182.600 73.100 ;
        RECT 183.800 70.800 184.200 72.100 ;
        RECT 185.400 70.800 185.800 73.100 ;
        RECT 188.100 70.800 188.600 72.100 ;
        RECT 189.800 70.800 190.200 72.100 ;
        RECT 192.600 70.800 193.000 73.000 ;
        RECT 0.200 70.200 195.800 70.800 ;
        RECT 1.400 67.900 1.800 70.200 ;
        RECT 3.000 67.900 3.400 70.200 ;
        RECT 4.600 67.900 5.000 70.200 ;
        RECT 6.200 67.900 6.600 70.200 ;
        RECT 7.800 67.900 8.200 70.200 ;
        RECT 9.400 67.900 9.800 70.200 ;
        RECT 11.000 68.000 11.400 70.200 ;
        RECT 13.800 68.900 14.200 70.200 ;
        RECT 15.400 68.900 15.900 70.200 ;
        RECT 18.200 67.900 18.600 70.200 ;
        RECT 21.400 68.300 21.800 70.200 ;
        RECT 23.800 68.900 24.200 70.200 ;
        RECT 25.400 67.900 25.800 70.200 ;
        RECT 28.100 68.900 28.600 70.200 ;
        RECT 29.800 68.900 30.200 70.200 ;
        RECT 32.600 68.000 33.000 70.200 ;
        RECT 35.800 68.300 36.200 70.200 ;
        RECT 38.200 68.900 38.600 70.200 ;
        RECT 39.800 67.900 40.200 70.200 ;
        RECT 42.500 68.900 43.000 70.200 ;
        RECT 44.200 68.900 44.600 70.200 ;
        RECT 47.000 68.000 47.400 70.200 ;
        RECT 50.200 68.900 50.600 70.200 ;
        RECT 53.400 67.900 53.800 70.200 ;
        RECT 54.500 67.900 54.900 70.200 ;
        RECT 56.600 68.900 57.000 70.200 ;
        RECT 59.000 68.300 59.400 70.200 ;
        RECT 60.600 68.900 61.000 70.200 ;
        RECT 62.200 68.900 62.600 70.200 ;
        RECT 63.800 68.000 64.200 70.200 ;
        RECT 66.600 68.900 67.000 70.200 ;
        RECT 68.200 68.900 68.700 70.200 ;
        RECT 71.000 67.900 71.400 70.200 ;
        RECT 73.400 67.700 73.800 70.200 ;
        RECT 76.000 67.500 76.400 70.200 ;
        RECT 78.200 68.000 78.600 70.200 ;
        RECT 81.000 68.900 81.400 70.200 ;
        RECT 82.600 68.900 83.100 70.200 ;
        RECT 85.400 67.900 85.800 70.200 ;
        RECT 87.000 68.900 87.400 70.200 ;
        RECT 88.600 68.900 89.000 70.200 ;
        RECT 90.200 67.900 90.600 70.200 ;
        RECT 92.900 68.900 93.400 70.200 ;
        RECT 94.600 68.900 95.000 70.200 ;
        RECT 97.400 68.000 97.800 70.200 ;
        RECT 101.400 68.000 101.800 70.200 ;
        RECT 104.200 68.900 104.600 70.200 ;
        RECT 105.800 68.900 106.300 70.200 ;
        RECT 108.600 67.900 109.000 70.200 ;
        RECT 110.200 68.900 110.600 70.200 ;
        RECT 111.800 68.900 112.200 70.200 ;
        RECT 113.400 68.900 113.800 70.200 ;
        RECT 115.000 67.900 115.400 70.200 ;
        RECT 117.700 68.900 118.200 70.200 ;
        RECT 119.400 68.900 119.800 70.200 ;
        RECT 122.200 68.000 122.600 70.200 ;
        RECT 123.800 67.900 124.200 70.200 ;
        RECT 125.400 67.900 125.800 70.200 ;
        RECT 127.000 67.900 127.400 70.200 ;
        RECT 128.600 67.900 129.000 70.200 ;
        RECT 130.200 67.900 130.600 70.200 ;
        RECT 131.800 67.900 132.200 70.200 ;
        RECT 134.500 68.900 135.000 70.200 ;
        RECT 136.200 68.900 136.600 70.200 ;
        RECT 139.000 68.000 139.400 70.200 ;
        RECT 140.600 67.900 141.000 70.200 ;
        RECT 142.200 67.900 142.600 70.200 ;
        RECT 143.800 67.900 144.200 70.200 ;
        RECT 145.400 67.900 145.800 70.200 ;
        RECT 147.000 67.900 147.400 70.200 ;
        RECT 150.200 67.900 150.600 70.200 ;
        RECT 152.900 68.000 153.300 70.200 ;
        RECT 155.800 67.900 156.200 70.200 ;
        RECT 158.500 68.000 158.900 70.200 ;
        RECT 162.200 67.900 162.600 70.200 ;
        RECT 165.400 66.900 165.800 70.200 ;
        RECT 166.200 67.900 166.600 70.200 ;
        RECT 167.800 67.900 168.200 70.200 ;
        RECT 170.200 67.900 170.600 70.200 ;
        RECT 171.800 68.900 172.200 70.200 ;
        RECT 173.400 68.900 173.800 70.200 ;
        RECT 175.800 68.300 176.200 70.200 ;
        RECT 177.400 68.900 177.800 70.200 ;
        RECT 179.000 68.900 179.400 70.200 ;
        RECT 180.600 67.900 181.000 70.200 ;
        RECT 183.300 68.900 183.800 70.200 ;
        RECT 185.000 68.900 185.400 70.200 ;
        RECT 187.800 68.000 188.200 70.200 ;
        RECT 190.200 67.900 190.600 70.200 ;
        RECT 192.600 67.900 193.000 70.200 ;
        RECT 2.200 65.800 2.600 66.600 ;
        RECT 0.600 50.800 1.000 53.100 ;
        RECT 2.200 50.800 2.600 53.100 ;
        RECT 3.800 50.800 4.200 53.100 ;
        RECT 5.400 50.800 5.800 53.100 ;
        RECT 7.000 50.800 7.400 53.100 ;
        RECT 7.800 50.800 8.200 52.100 ;
        RECT 9.400 50.800 9.800 52.100 ;
        RECT 11.000 50.800 11.400 53.300 ;
        RECT 13.600 50.800 14.000 53.500 ;
        RECT 15.000 50.800 15.400 53.100 ;
        RECT 17.400 50.800 17.800 53.100 ;
        RECT 19.000 50.800 19.400 53.100 ;
        RECT 20.600 50.800 21.000 52.100 ;
        RECT 22.200 50.800 22.600 52.100 ;
        RECT 23.800 50.800 24.200 53.300 ;
        RECT 26.400 50.800 26.800 53.500 ;
        RECT 27.800 50.800 28.200 53.100 ;
        RECT 31.000 51.100 31.500 52.800 ;
        RECT 31.100 50.800 31.500 51.100 ;
        RECT 34.100 50.800 34.600 52.800 ;
        RECT 35.800 50.800 36.200 52.100 ;
        RECT 38.200 50.800 38.600 52.700 ;
        RECT 42.200 50.800 42.600 53.100 ;
        RECT 43.000 50.800 43.400 52.100 ;
        RECT 47.000 50.800 47.400 52.700 ;
        RECT 49.400 50.800 49.800 53.100 ;
        RECT 52.600 50.800 53.000 53.000 ;
        RECT 55.400 50.800 55.800 52.100 ;
        RECT 57.000 50.800 57.500 52.100 ;
        RECT 59.800 50.800 60.200 53.100 ;
        RECT 62.200 50.800 62.600 53.000 ;
        RECT 65.000 50.800 65.400 52.100 ;
        RECT 66.600 50.800 67.100 52.100 ;
        RECT 69.400 50.800 69.800 53.100 ;
        RECT 71.000 50.800 71.400 52.100 ;
        RECT 72.600 50.800 73.000 52.100 ;
        RECT 73.400 50.800 73.800 52.100 ;
        RECT 75.000 50.800 75.400 52.100 ;
        RECT 76.600 50.800 77.000 53.300 ;
        RECT 79.200 50.800 79.600 53.500 ;
        RECT 80.800 50.800 81.200 53.100 ;
        RECT 83.800 50.800 84.200 53.100 ;
        RECT 84.600 50.800 85.000 52.100 ;
        RECT 86.700 50.800 87.100 53.100 ;
        RECT 87.800 50.800 88.200 52.100 ;
        RECT 89.400 50.800 89.800 52.100 ;
        RECT 90.200 50.800 90.600 53.100 ;
        RECT 92.600 50.800 93.000 52.100 ;
        RECT 96.600 50.800 97.000 52.100 ;
        RECT 98.200 50.800 98.600 51.900 ;
        RECT 102.400 50.800 102.800 53.100 ;
        RECT 105.400 50.800 105.800 53.100 ;
        RECT 106.200 50.800 106.600 52.100 ;
        RECT 107.800 50.800 108.200 52.100 ;
        RECT 109.900 50.800 110.300 53.000 ;
        RECT 111.800 50.800 112.200 53.100 ;
        RECT 114.800 50.800 115.200 53.100 ;
        RECT 116.600 50.800 117.000 52.900 ;
        RECT 118.200 50.800 118.600 52.100 ;
        RECT 119.300 50.800 119.700 53.100 ;
        RECT 121.400 50.800 121.800 52.100 ;
        RECT 123.000 50.800 123.400 53.100 ;
        RECT 125.400 50.800 125.800 53.000 ;
        RECT 128.200 50.800 128.600 52.100 ;
        RECT 129.800 50.800 130.300 52.100 ;
        RECT 132.600 50.800 133.000 53.100 ;
        RECT 134.200 50.800 134.600 52.100 ;
        RECT 136.300 50.800 136.700 53.100 ;
        RECT 137.400 50.800 137.800 52.100 ;
        RECT 139.500 50.800 139.900 53.100 ;
        RECT 140.600 50.800 141.000 52.100 ;
        RECT 142.200 50.800 142.600 53.100 ;
        RECT 144.900 50.800 145.300 53.100 ;
        RECT 147.000 50.800 147.400 52.100 ;
        RECT 151.000 50.800 151.400 52.700 ;
        RECT 152.600 50.800 153.000 53.100 ;
        RECT 155.000 50.800 155.500 52.800 ;
        RECT 158.100 51.100 158.600 52.800 ;
        RECT 158.100 50.800 158.500 51.100 ;
        RECT 159.800 50.800 160.200 52.100 ;
        RECT 161.400 50.800 161.800 52.100 ;
        RECT 164.600 50.800 165.000 54.100 ;
        RECT 165.400 50.800 165.800 53.100 ;
        RECT 167.800 50.800 168.200 52.100 ;
        RECT 169.400 50.800 169.800 52.100 ;
        RECT 170.200 50.800 170.600 54.100 ;
        RECT 173.400 50.800 173.800 52.100 ;
        RECT 176.600 50.800 177.000 52.700 ;
        RECT 178.200 50.800 178.600 52.100 ;
        RECT 179.800 50.800 180.200 52.100 ;
        RECT 182.200 50.800 182.600 52.700 ;
        RECT 184.600 50.800 185.000 53.100 ;
        RECT 187.300 50.800 187.800 52.100 ;
        RECT 189.000 50.800 189.400 52.100 ;
        RECT 191.800 50.800 192.200 53.000 ;
        RECT 194.200 50.800 194.600 52.100 ;
        RECT 0.200 50.200 195.800 50.800 ;
        RECT 1.400 47.900 1.800 50.200 ;
        RECT 3.800 48.000 4.200 50.200 ;
        RECT 6.600 48.900 7.000 50.200 ;
        RECT 8.200 48.900 8.700 50.200 ;
        RECT 11.000 47.900 11.400 50.200 ;
        RECT 12.600 48.900 13.000 50.200 ;
        RECT 14.200 48.900 14.600 50.200 ;
        RECT 15.800 47.900 16.200 50.200 ;
        RECT 18.500 48.900 19.000 50.200 ;
        RECT 20.200 48.900 20.600 50.200 ;
        RECT 23.000 48.000 23.400 50.200 ;
        RECT 25.400 47.900 25.800 50.200 ;
        RECT 28.100 48.900 28.600 50.200 ;
        RECT 29.800 48.900 30.200 50.200 ;
        RECT 32.600 48.000 33.000 50.200 ;
        RECT 37.400 49.100 37.800 50.200 ;
        RECT 39.000 48.900 39.400 50.200 ;
        RECT 41.400 48.200 41.900 50.200 ;
        RECT 44.500 49.900 44.900 50.200 ;
        RECT 44.500 48.200 45.000 49.900 ;
        RECT 48.600 48.000 49.000 50.200 ;
        RECT 51.400 48.900 51.800 50.200 ;
        RECT 53.000 48.900 53.500 50.200 ;
        RECT 55.800 47.900 56.200 50.200 ;
        RECT 57.400 47.900 57.800 50.200 ;
        RECT 59.000 47.900 59.400 50.200 ;
        RECT 60.600 47.900 61.000 50.200 ;
        RECT 62.200 47.900 62.600 50.200 ;
        RECT 63.800 47.900 64.200 50.200 ;
        RECT 65.400 47.900 65.800 50.200 ;
        RECT 67.800 48.900 68.200 50.200 ;
        RECT 69.400 48.000 69.800 50.200 ;
        RECT 72.200 48.900 72.600 50.200 ;
        RECT 73.800 48.900 74.300 50.200 ;
        RECT 76.600 47.900 77.000 50.200 ;
        RECT 79.800 48.300 80.200 50.200 ;
        RECT 81.400 47.900 81.800 50.200 ;
        RECT 83.800 48.900 84.200 50.200 ;
        RECT 85.400 48.900 85.800 50.200 ;
        RECT 87.000 47.900 87.400 50.200 ;
        RECT 87.800 48.900 88.200 50.200 ;
        RECT 89.400 48.900 89.800 50.200 ;
        RECT 90.200 47.900 90.600 50.200 ;
        RECT 92.600 47.900 93.000 50.200 ;
        RECT 99.000 49.100 99.400 50.200 ;
        RECT 100.600 48.900 101.000 50.200 ;
        RECT 103.000 48.900 103.400 50.200 ;
        RECT 104.600 47.900 105.000 50.200 ;
        RECT 107.000 48.900 107.400 50.200 ;
        RECT 108.600 49.100 109.000 50.200 ;
        RECT 112.800 47.900 113.200 50.200 ;
        RECT 115.800 47.900 116.200 50.200 ;
        RECT 116.900 47.900 117.300 50.200 ;
        RECT 119.000 48.900 119.400 50.200 ;
        RECT 120.600 48.000 121.000 50.200 ;
        RECT 123.400 48.900 123.800 50.200 ;
        RECT 125.000 48.900 125.500 50.200 ;
        RECT 127.800 47.900 128.200 50.200 ;
        RECT 130.200 47.900 130.600 50.200 ;
        RECT 132.900 48.900 133.400 50.200 ;
        RECT 134.600 48.900 135.000 50.200 ;
        RECT 137.400 48.000 137.800 50.200 ;
        RECT 139.800 48.000 140.200 50.200 ;
        RECT 142.600 48.900 143.000 50.200 ;
        RECT 144.200 48.900 144.700 50.200 ;
        RECT 147.000 47.900 147.400 50.200 ;
        RECT 150.200 48.900 150.600 50.200 ;
        RECT 151.800 48.900 152.200 50.200 ;
        RECT 152.600 48.900 153.000 50.200 ;
        RECT 154.200 48.900 154.600 50.200 ;
        RECT 157.400 46.900 157.800 50.200 ;
        RECT 159.000 48.000 159.400 50.200 ;
        RECT 161.800 48.900 162.200 50.200 ;
        RECT 163.400 48.900 163.900 50.200 ;
        RECT 166.200 47.900 166.600 50.200 ;
        RECT 169.400 47.900 169.800 50.200 ;
        RECT 170.200 48.900 170.600 50.200 ;
        RECT 171.800 48.900 172.200 50.200 ;
        RECT 173.400 47.900 173.800 50.200 ;
        RECT 176.100 48.900 176.600 50.200 ;
        RECT 177.800 48.900 178.200 50.200 ;
        RECT 180.600 48.000 181.000 50.200 ;
        RECT 183.000 47.900 183.400 50.200 ;
        RECT 185.700 48.900 186.200 50.200 ;
        RECT 187.400 48.900 187.800 50.200 ;
        RECT 190.200 48.000 190.600 50.200 ;
        RECT 192.600 47.900 193.000 50.200 ;
        RECT 2.200 45.800 2.600 46.600 ;
        RECT 191.800 45.800 192.200 46.600 ;
        RECT 191.800 34.400 192.200 35.200 ;
        RECT 1.400 30.800 1.800 33.000 ;
        RECT 4.200 30.800 4.600 32.100 ;
        RECT 5.800 30.800 6.300 32.100 ;
        RECT 8.600 30.800 9.000 33.100 ;
        RECT 11.000 30.800 11.400 33.000 ;
        RECT 13.800 30.800 14.200 32.100 ;
        RECT 15.400 30.800 15.900 32.100 ;
        RECT 18.200 30.800 18.600 33.100 ;
        RECT 20.600 30.800 21.000 33.100 ;
        RECT 23.300 30.800 23.800 32.100 ;
        RECT 25.000 30.800 25.400 32.100 ;
        RECT 27.800 30.800 28.200 33.000 ;
        RECT 30.200 30.800 30.600 33.000 ;
        RECT 33.000 30.800 33.400 32.100 ;
        RECT 34.600 30.800 35.100 32.100 ;
        RECT 37.400 30.800 37.800 33.100 ;
        RECT 40.300 30.800 40.700 33.000 ;
        RECT 43.000 30.800 43.400 32.700 ;
        RECT 48.900 30.800 49.300 33.000 ;
        RECT 51.000 30.800 51.400 32.100 ;
        RECT 52.600 30.800 53.000 32.100 ;
        RECT 54.200 30.800 54.600 33.000 ;
        RECT 57.000 30.800 57.400 32.100 ;
        RECT 58.600 30.800 59.100 32.100 ;
        RECT 61.400 30.800 61.800 33.100 ;
        RECT 63.800 30.800 64.200 32.900 ;
        RECT 65.400 30.800 65.800 32.100 ;
        RECT 66.200 30.800 66.600 32.100 ;
        RECT 67.800 30.800 68.200 32.100 ;
        RECT 69.400 30.800 69.800 32.100 ;
        RECT 71.800 30.800 72.200 33.100 ;
        RECT 73.700 30.800 74.100 33.000 ;
        RECT 75.800 30.800 76.200 32.100 ;
        RECT 77.400 30.800 77.800 32.100 ;
        RECT 78.200 30.800 78.600 32.100 ;
        RECT 80.600 30.800 81.000 33.100 ;
        RECT 83.300 30.800 83.800 32.100 ;
        RECT 85.000 30.800 85.400 32.100 ;
        RECT 87.800 30.800 88.200 33.000 ;
        RECT 90.200 30.800 90.600 33.100 ;
        RECT 92.900 30.800 93.400 32.100 ;
        RECT 94.600 30.800 95.000 32.100 ;
        RECT 97.400 30.800 97.800 33.000 ;
        RECT 101.700 30.800 102.100 33.000 ;
        RECT 104.600 30.800 105.000 32.100 ;
        RECT 106.200 30.800 106.600 31.900 ;
        RECT 110.200 30.800 110.600 32.100 ;
        RECT 111.800 30.800 112.200 32.100 ;
        RECT 113.400 30.800 113.800 33.000 ;
        RECT 116.200 30.800 116.600 32.100 ;
        RECT 117.800 30.800 118.300 32.100 ;
        RECT 120.600 30.800 121.000 33.100 ;
        RECT 122.200 30.800 122.600 32.100 ;
        RECT 123.800 30.800 124.200 32.100 ;
        RECT 125.400 30.800 125.800 33.000 ;
        RECT 128.200 30.800 128.600 32.100 ;
        RECT 129.800 30.800 130.300 32.100 ;
        RECT 132.600 30.800 133.000 33.100 ;
        RECT 135.000 30.800 135.400 33.100 ;
        RECT 137.400 30.800 137.800 33.100 ;
        RECT 139.000 30.800 139.400 33.100 ;
        RECT 140.600 30.800 141.000 33.100 ;
        RECT 142.200 30.800 142.600 33.100 ;
        RECT 143.800 30.800 144.200 33.100 ;
        RECT 145.400 30.800 145.800 33.100 ;
        RECT 148.600 30.800 149.000 33.100 ;
        RECT 151.300 30.800 151.800 32.100 ;
        RECT 153.000 30.800 153.400 32.100 ;
        RECT 155.800 30.800 156.200 33.000 ;
        RECT 158.200 30.800 158.600 33.100 ;
        RECT 160.900 30.800 161.400 32.100 ;
        RECT 162.600 30.800 163.000 32.100 ;
        RECT 165.400 30.800 165.800 33.000 ;
        RECT 167.000 30.800 167.400 32.100 ;
        RECT 169.100 30.800 169.500 33.100 ;
        RECT 171.000 30.800 171.400 33.000 ;
        RECT 173.800 30.800 174.200 32.100 ;
        RECT 175.400 30.800 175.900 32.100 ;
        RECT 178.200 30.800 178.600 33.100 ;
        RECT 180.600 30.800 181.000 33.100 ;
        RECT 183.300 30.800 183.800 32.100 ;
        RECT 185.000 30.800 185.400 32.100 ;
        RECT 187.800 30.800 188.200 33.000 ;
        RECT 190.200 30.800 190.600 33.100 ;
        RECT 192.600 30.800 193.000 33.100 ;
        RECT 0.200 30.200 195.800 30.800 ;
        RECT 0.600 28.900 1.000 30.200 ;
        RECT 2.200 28.100 2.600 30.200 ;
        RECT 3.800 28.900 4.200 30.200 ;
        RECT 5.400 28.100 5.800 30.200 ;
        RECT 7.000 28.900 7.400 30.200 ;
        RECT 9.400 27.900 9.800 30.200 ;
        RECT 12.100 28.900 12.600 30.200 ;
        RECT 13.800 28.900 14.200 30.200 ;
        RECT 16.600 28.000 17.000 30.200 ;
        RECT 19.000 27.900 19.400 30.200 ;
        RECT 21.700 28.900 22.200 30.200 ;
        RECT 23.400 28.900 23.800 30.200 ;
        RECT 26.200 28.000 26.600 30.200 ;
        RECT 28.600 27.900 29.000 30.200 ;
        RECT 31.300 28.900 31.800 30.200 ;
        RECT 33.000 28.900 33.400 30.200 ;
        RECT 35.800 28.000 36.200 30.200 ;
        RECT 37.400 28.900 37.800 30.200 ;
        RECT 39.000 28.900 39.400 30.200 ;
        RECT 40.600 27.900 41.000 30.200 ;
        RECT 43.300 28.900 43.800 30.200 ;
        RECT 45.000 28.900 45.400 30.200 ;
        RECT 47.800 28.000 48.200 30.200 ;
        RECT 52.300 28.000 52.700 30.200 ;
        RECT 55.000 28.000 55.400 30.200 ;
        RECT 57.800 28.900 58.200 30.200 ;
        RECT 59.400 28.900 59.900 30.200 ;
        RECT 62.200 27.900 62.600 30.200 ;
        RECT 64.600 27.900 65.000 30.200 ;
        RECT 67.000 28.100 67.400 30.200 ;
        RECT 68.600 28.900 69.000 30.200 ;
        RECT 69.400 28.900 69.800 30.200 ;
        RECT 71.000 28.900 71.400 30.200 ;
        RECT 71.800 28.900 72.200 30.200 ;
        RECT 73.400 26.900 73.800 30.200 ;
        RECT 76.600 27.900 77.000 30.200 ;
        RECT 79.000 28.000 79.400 30.200 ;
        RECT 81.800 28.900 82.200 30.200 ;
        RECT 83.400 28.900 83.900 30.200 ;
        RECT 86.200 27.900 86.600 30.200 ;
        RECT 88.600 28.000 89.000 30.200 ;
        RECT 91.400 28.900 91.800 30.200 ;
        RECT 93.000 28.900 93.500 30.200 ;
        RECT 95.800 27.900 96.200 30.200 ;
        RECT 100.300 28.000 100.700 30.200 ;
        RECT 103.000 28.000 103.400 30.200 ;
        RECT 105.800 28.900 106.200 30.200 ;
        RECT 107.400 28.900 107.900 30.200 ;
        RECT 110.200 27.900 110.600 30.200 ;
        RECT 112.600 28.000 113.000 30.200 ;
        RECT 115.400 28.900 115.800 30.200 ;
        RECT 117.000 28.900 117.500 30.200 ;
        RECT 119.800 27.900 120.200 30.200 ;
        RECT 121.400 28.900 121.800 30.200 ;
        RECT 123.000 27.900 123.400 30.200 ;
        RECT 124.600 27.900 125.000 30.200 ;
        RECT 126.200 27.900 126.600 30.200 ;
        RECT 127.800 27.900 128.200 30.200 ;
        RECT 129.400 27.900 129.800 30.200 ;
        RECT 130.200 28.900 130.600 30.200 ;
        RECT 131.800 28.900 132.200 30.200 ;
        RECT 133.400 28.900 133.800 30.200 ;
        RECT 135.000 27.900 135.400 30.200 ;
        RECT 137.700 28.900 138.200 30.200 ;
        RECT 139.400 28.900 139.800 30.200 ;
        RECT 142.200 28.000 142.600 30.200 ;
        RECT 146.200 27.900 146.600 30.200 ;
        RECT 148.900 28.900 149.400 30.200 ;
        RECT 150.600 28.900 151.000 30.200 ;
        RECT 153.400 28.000 153.800 30.200 ;
        RECT 155.800 27.900 156.200 30.200 ;
        RECT 158.500 28.900 159.000 30.200 ;
        RECT 160.200 28.900 160.600 30.200 ;
        RECT 163.000 28.000 163.400 30.200 ;
        RECT 166.200 28.300 166.600 30.200 ;
        RECT 168.600 28.000 169.000 30.200 ;
        RECT 171.400 28.900 171.800 30.200 ;
        RECT 173.000 28.900 173.500 30.200 ;
        RECT 175.800 27.900 176.200 30.200 ;
        RECT 177.400 28.900 177.800 30.200 ;
        RECT 179.000 28.900 179.400 30.200 ;
        RECT 180.600 27.900 181.000 30.200 ;
        RECT 183.300 28.900 183.800 30.200 ;
        RECT 185.000 28.900 185.400 30.200 ;
        RECT 187.800 28.000 188.200 30.200 ;
        RECT 190.200 27.900 190.600 30.200 ;
        RECT 192.600 27.900 193.000 30.200 ;
        RECT 191.000 25.800 191.400 26.600 ;
        RECT 2.200 14.400 2.600 15.200 ;
        RECT 94.200 14.400 94.600 15.200 ;
        RECT 1.400 10.800 1.800 13.100 ;
        RECT 3.800 10.800 4.200 13.000 ;
        RECT 6.600 10.800 7.000 12.100 ;
        RECT 8.200 10.800 8.700 12.100 ;
        RECT 11.000 10.800 11.400 13.100 ;
        RECT 12.600 10.800 13.000 12.100 ;
        RECT 14.200 10.800 14.600 12.100 ;
        RECT 15.800 10.800 16.200 13.100 ;
        RECT 18.500 10.800 19.000 12.100 ;
        RECT 20.200 10.800 20.600 12.100 ;
        RECT 23.000 10.800 23.400 13.000 ;
        RECT 24.600 10.800 25.000 12.100 ;
        RECT 26.200 10.800 26.600 12.100 ;
        RECT 27.300 10.800 27.700 13.100 ;
        RECT 29.400 10.800 29.800 12.100 ;
        RECT 30.200 10.800 30.600 13.100 ;
        RECT 32.600 10.800 33.000 12.100 ;
        RECT 34.200 10.800 34.600 12.100 ;
        RECT 35.800 10.800 36.200 13.000 ;
        RECT 38.600 10.800 39.000 12.100 ;
        RECT 40.200 10.800 40.700 12.100 ;
        RECT 43.000 10.800 43.400 13.100 ;
        RECT 47.500 10.800 47.900 13.000 ;
        RECT 50.200 10.800 50.600 13.000 ;
        RECT 53.000 10.800 53.400 12.100 ;
        RECT 54.600 10.800 55.100 12.100 ;
        RECT 57.400 10.800 57.800 13.100 ;
        RECT 59.000 10.800 59.400 13.100 ;
        RECT 60.600 10.800 61.000 13.100 ;
        RECT 62.200 10.800 62.600 13.100 ;
        RECT 63.800 10.800 64.200 13.100 ;
        RECT 65.400 10.800 65.800 13.100 ;
        RECT 67.000 10.800 67.400 13.100 ;
        RECT 69.700 10.800 70.200 12.100 ;
        RECT 71.400 10.800 71.800 12.100 ;
        RECT 74.200 10.800 74.600 13.000 ;
        RECT 76.900 10.800 77.300 13.000 ;
        RECT 80.600 10.800 81.000 13.100 ;
        RECT 81.400 10.800 81.800 12.100 ;
        RECT 83.000 10.800 83.400 12.100 ;
        RECT 83.800 10.800 84.200 12.100 ;
        RECT 85.700 10.800 86.100 13.100 ;
        RECT 87.800 10.800 88.200 12.100 ;
        RECT 90.200 10.800 90.600 12.700 ;
        RECT 91.800 10.800 92.200 12.100 ;
        RECT 93.400 10.800 93.800 12.100 ;
        RECT 95.000 10.800 95.400 13.100 ;
        RECT 99.000 10.800 99.400 12.100 ;
        RECT 100.600 10.800 101.000 11.900 ;
        RECT 104.600 10.800 105.000 13.100 ;
        RECT 107.800 10.800 108.200 12.700 ;
        RECT 110.200 10.800 110.600 12.100 ;
        RECT 111.800 10.800 112.200 12.100 ;
        RECT 112.600 10.800 113.000 12.100 ;
        RECT 114.700 10.800 115.100 13.100 ;
        RECT 116.600 10.800 117.000 13.100 ;
        RECT 117.400 10.800 117.800 12.100 ;
        RECT 119.000 10.800 119.400 12.100 ;
        RECT 120.600 10.800 121.000 12.100 ;
        RECT 122.200 10.800 122.600 13.000 ;
        RECT 125.000 10.800 125.400 12.100 ;
        RECT 126.600 10.800 127.100 12.100 ;
        RECT 129.400 10.800 129.800 13.100 ;
        RECT 131.000 10.800 131.400 12.100 ;
        RECT 132.600 10.800 133.000 12.100 ;
        RECT 135.000 10.800 135.400 12.700 ;
        RECT 137.400 10.800 137.800 12.700 ;
        RECT 140.100 10.800 140.500 13.100 ;
        RECT 142.200 10.800 142.600 12.100 ;
        RECT 143.800 10.800 144.200 13.100 ;
        RECT 146.500 10.800 147.000 12.100 ;
        RECT 148.200 10.800 148.600 12.100 ;
        RECT 151.000 10.800 151.400 13.000 ;
        RECT 154.200 10.800 154.600 13.100 ;
        RECT 156.600 10.800 157.000 12.900 ;
        RECT 158.200 10.800 158.600 12.100 ;
        RECT 159.800 10.800 160.200 13.100 ;
        RECT 162.500 10.800 163.000 12.100 ;
        RECT 164.200 10.800 164.600 12.100 ;
        RECT 167.000 10.800 167.400 13.000 ;
        RECT 170.200 10.800 170.600 13.100 ;
        RECT 171.000 10.800 171.400 12.100 ;
        RECT 173.100 10.800 173.500 13.100 ;
        RECT 175.000 10.800 175.400 13.100 ;
        RECT 177.400 10.800 177.800 13.100 ;
        RECT 179.800 10.800 180.200 12.700 ;
        RECT 181.400 10.800 181.800 12.100 ;
        RECT 183.000 10.800 183.400 12.100 ;
        RECT 183.800 10.800 184.200 12.100 ;
        RECT 186.200 10.800 186.600 13.100 ;
        RECT 188.900 10.800 189.400 12.100 ;
        RECT 190.600 10.800 191.000 12.100 ;
        RECT 193.400 10.800 193.800 13.000 ;
        RECT 0.200 10.200 195.800 10.800 ;
        RECT 0.600 8.900 1.000 10.200 ;
        RECT 3.000 8.300 3.400 10.200 ;
        RECT 5.400 8.900 5.800 10.200 ;
        RECT 7.000 8.900 7.400 10.200 ;
        RECT 11.000 9.100 11.400 10.200 ;
        RECT 12.600 8.900 13.000 10.200 ;
        RECT 14.200 8.900 14.600 10.200 ;
        RECT 15.800 8.900 16.200 10.200 ;
        RECT 18.200 7.900 18.600 10.200 ;
        RECT 20.600 8.300 21.000 10.200 ;
        RECT 22.200 7.900 22.600 10.200 ;
        RECT 23.800 8.900 24.200 10.200 ;
        RECT 25.400 8.900 25.800 10.200 ;
        RECT 29.400 9.100 29.800 10.200 ;
        RECT 31.000 8.900 31.400 10.200 ;
        RECT 34.200 7.900 34.600 10.200 ;
        RECT 35.800 8.000 36.200 10.200 ;
        RECT 38.600 8.900 39.000 10.200 ;
        RECT 40.200 8.900 40.700 10.200 ;
        RECT 43.000 7.900 43.400 10.200 ;
        RECT 47.000 8.300 47.400 10.200 ;
        RECT 49.400 8.900 49.800 10.200 ;
        RECT 51.000 8.900 51.400 10.200 ;
        RECT 51.800 8.900 52.200 10.200 ;
        RECT 54.200 8.300 54.600 10.200 ;
        RECT 57.400 7.900 57.800 10.200 ;
        RECT 59.300 7.900 59.700 10.200 ;
        RECT 61.400 8.900 61.800 10.200 ;
        RECT 62.200 7.900 62.600 10.200 ;
        RECT 65.400 7.900 65.800 10.200 ;
        RECT 68.100 8.900 68.600 10.200 ;
        RECT 69.800 8.900 70.200 10.200 ;
        RECT 72.600 8.000 73.000 10.200 ;
        RECT 74.200 8.900 74.600 10.200 ;
        RECT 76.100 7.900 76.500 10.200 ;
        RECT 78.200 8.900 78.600 10.200 ;
        RECT 79.000 8.900 79.400 10.200 ;
        RECT 80.600 8.100 81.000 10.200 ;
        RECT 82.200 8.900 82.600 10.200 ;
        RECT 83.800 6.900 84.200 10.200 ;
        RECT 88.600 7.900 89.000 10.200 ;
        RECT 90.200 7.900 90.600 10.200 ;
        RECT 92.900 8.900 93.400 10.200 ;
        RECT 94.600 8.900 95.000 10.200 ;
        RECT 97.400 8.000 97.800 10.200 ;
        RECT 100.600 8.900 101.000 10.200 ;
        RECT 102.200 8.900 102.600 10.200 ;
        RECT 104.600 7.900 105.000 10.200 ;
        RECT 106.500 8.000 106.900 10.200 ;
        RECT 109.400 8.000 109.800 10.200 ;
        RECT 112.200 8.900 112.600 10.200 ;
        RECT 113.800 8.900 114.300 10.200 ;
        RECT 116.600 7.900 117.000 10.200 ;
        RECT 119.800 7.900 120.200 10.200 ;
        RECT 120.600 8.900 121.000 10.200 ;
        RECT 122.200 8.900 122.600 10.200 ;
        RECT 123.800 8.300 124.200 10.200 ;
        RECT 126.200 7.900 126.600 10.200 ;
        RECT 129.400 7.900 129.800 10.200 ;
        RECT 132.100 8.900 132.600 10.200 ;
        RECT 133.800 8.900 134.200 10.200 ;
        RECT 136.600 8.000 137.000 10.200 ;
        RECT 139.500 8.000 139.900 10.200 ;
        RECT 142.200 7.900 142.600 10.200 ;
        RECT 144.900 8.900 145.400 10.200 ;
        RECT 146.600 8.900 147.000 10.200 ;
        RECT 149.400 8.000 149.800 10.200 ;
        RECT 153.400 8.000 153.800 10.200 ;
        RECT 156.200 8.900 156.600 10.200 ;
        RECT 157.800 8.900 158.300 10.200 ;
        RECT 160.600 7.900 161.000 10.200 ;
        RECT 162.200 8.900 162.600 10.200 ;
        RECT 163.800 8.900 164.200 10.200 ;
        RECT 165.400 7.900 165.800 10.200 ;
        RECT 167.800 8.300 168.200 10.200 ;
        RECT 170.200 8.900 170.600 10.200 ;
        RECT 171.800 8.900 172.200 10.200 ;
        RECT 173.400 8.000 173.800 10.200 ;
        RECT 176.200 8.900 176.600 10.200 ;
        RECT 177.800 8.900 178.300 10.200 ;
        RECT 180.600 7.900 181.000 10.200 ;
        RECT 182.200 8.900 182.600 10.200 ;
        RECT 183.800 8.900 184.200 10.200 ;
        RECT 185.400 7.900 185.800 10.200 ;
        RECT 188.100 8.900 188.600 10.200 ;
        RECT 189.800 8.900 190.200 10.200 ;
        RECT 192.600 8.000 193.000 10.200 ;
        RECT 56.600 5.800 57.000 6.600 ;
        RECT 164.600 5.800 165.000 6.600 ;
      LAYER via1 ;
        RECT 97.000 170.300 97.400 170.700 ;
        RECT 97.700 170.300 98.100 170.700 ;
        RECT 97.000 150.300 97.400 150.700 ;
        RECT 97.700 150.300 98.100 150.700 ;
        RECT 27.000 134.800 27.400 135.200 ;
        RECT 189.400 134.800 189.800 135.200 ;
        RECT 27.800 132.700 28.200 133.100 ;
        RECT 190.200 132.700 190.600 133.100 ;
        RECT 97.000 130.300 97.400 130.700 ;
        RECT 97.700 130.300 98.100 130.700 ;
        RECT 191.800 114.800 192.200 115.200 ;
        RECT 97.000 110.300 97.400 110.700 ;
        RECT 97.700 110.300 98.100 110.700 ;
        RECT 191.800 109.800 192.200 110.200 ;
        RECT 192.600 94.800 193.000 95.200 ;
        RECT 97.000 90.300 97.400 90.700 ;
        RECT 97.700 90.300 98.100 90.700 ;
        RECT 192.600 89.800 193.000 90.200 ;
        RECT 97.000 70.300 97.400 70.700 ;
        RECT 97.700 70.300 98.100 70.700 ;
        RECT 97.000 50.300 97.400 50.700 ;
        RECT 97.700 50.300 98.100 50.700 ;
        RECT 191.800 34.800 192.200 35.200 ;
        RECT 192.600 32.700 193.000 33.100 ;
        RECT 97.000 30.300 97.400 30.700 ;
        RECT 97.700 30.300 98.100 30.700 ;
        RECT 2.200 14.800 2.600 15.200 ;
        RECT 94.200 14.800 94.600 15.200 ;
        RECT 1.400 12.700 1.800 13.100 ;
        RECT 95.000 12.700 95.400 13.100 ;
        RECT 97.000 10.300 97.400 10.700 ;
        RECT 97.700 10.300 98.100 10.700 ;
      LAYER metal2 ;
        RECT 96.800 170.300 98.400 170.700 ;
        RECT 105.400 168.100 105.800 168.300 ;
        RECT 104.600 167.900 105.800 168.100 ;
        RECT 186.200 168.100 186.600 168.300 ;
        RECT 104.600 167.800 105.700 167.900 ;
        RECT 186.200 167.800 187.300 168.100 ;
        RECT 104.600 166.200 104.900 167.800 ;
        RECT 187.000 166.200 187.300 167.800 ;
        RECT 104.600 165.800 105.000 166.200 ;
        RECT 187.000 165.800 187.400 166.200 ;
        RECT 96.800 150.300 98.400 150.700 ;
        RECT 27.000 134.800 27.400 135.200 ;
        RECT 189.400 134.800 189.800 135.200 ;
        RECT 27.000 133.100 27.300 134.800 ;
        RECT 189.400 133.100 189.700 134.800 ;
        RECT 27.000 132.800 28.200 133.100 ;
        RECT 189.400 132.800 190.600 133.100 ;
        RECT 27.800 132.700 28.200 132.800 ;
        RECT 190.200 132.700 190.600 132.800 ;
        RECT 96.800 130.300 98.400 130.700 ;
        RECT 191.800 114.800 192.200 115.200 ;
        RECT 96.800 110.300 98.400 110.700 ;
        RECT 191.800 110.200 192.100 114.800 ;
        RECT 191.800 109.800 192.200 110.200 ;
        RECT 192.600 94.800 193.000 95.200 ;
        RECT 155.000 90.800 155.400 91.200 ;
        RECT 96.800 90.300 98.400 90.700 ;
        RECT 155.000 86.200 155.300 90.800 ;
        RECT 192.600 90.200 192.900 94.800 ;
        RECT 192.600 89.800 193.000 90.200 ;
        RECT 190.200 88.100 190.600 88.300 ;
        RECT 189.400 87.900 190.600 88.100 ;
        RECT 189.400 87.800 190.500 87.900 ;
        RECT 189.400 86.200 189.700 87.800 ;
        RECT 155.000 85.800 155.400 86.200 ;
        RECT 189.400 85.800 189.800 86.200 ;
        RECT 2.200 70.800 2.600 71.200 ;
        RECT 2.200 66.200 2.500 70.800 ;
        RECT 96.800 70.300 98.400 70.700 ;
        RECT 2.200 65.800 2.600 66.200 ;
        RECT 2.200 50.800 2.600 51.200 ;
        RECT 191.800 50.800 192.200 51.200 ;
        RECT 2.200 46.200 2.500 50.800 ;
        RECT 96.800 50.300 98.400 50.700 ;
        RECT 191.800 46.200 192.100 50.800 ;
        RECT 2.200 45.800 2.600 46.200 ;
        RECT 191.800 45.800 192.200 46.200 ;
        RECT 191.800 34.800 192.200 35.200 ;
        RECT 191.800 33.100 192.100 34.800 ;
        RECT 191.800 32.800 193.000 33.100 ;
        RECT 192.600 32.700 193.000 32.800 ;
        RECT 96.800 30.300 98.400 30.700 ;
        RECT 190.200 28.100 190.600 28.300 ;
        RECT 190.200 27.800 191.300 28.100 ;
        RECT 191.000 26.200 191.300 27.800 ;
        RECT 191.000 25.800 191.400 26.200 ;
        RECT 2.200 14.800 2.600 15.200 ;
        RECT 94.200 14.800 94.600 15.200 ;
        RECT 2.200 13.100 2.500 14.800 ;
        RECT 1.400 12.800 2.500 13.100 ;
        RECT 94.200 13.100 94.500 14.800 ;
        RECT 94.200 12.800 95.400 13.100 ;
        RECT 1.400 12.700 1.800 12.800 ;
        RECT 95.000 12.700 95.400 12.800 ;
        RECT 96.800 10.300 98.400 10.700 ;
        RECT 57.400 8.100 57.800 8.300 ;
        RECT 165.400 8.100 165.800 8.300 ;
        RECT 56.600 7.900 57.800 8.100 ;
        RECT 164.600 7.900 165.800 8.100 ;
        RECT 56.600 7.800 57.700 7.900 ;
        RECT 164.600 7.800 165.700 7.900 ;
        RECT 56.600 6.200 56.900 7.800 ;
        RECT 164.600 6.200 164.900 7.800 ;
        RECT 56.600 5.800 57.000 6.200 ;
        RECT 164.600 5.800 165.000 6.200 ;
      LAYER via2 ;
        RECT 97.000 170.300 97.400 170.700 ;
        RECT 97.700 170.300 98.100 170.700 ;
        RECT 97.000 150.300 97.400 150.700 ;
        RECT 97.700 150.300 98.100 150.700 ;
        RECT 97.000 130.300 97.400 130.700 ;
        RECT 97.700 130.300 98.100 130.700 ;
        RECT 97.000 110.300 97.400 110.700 ;
        RECT 97.700 110.300 98.100 110.700 ;
        RECT 97.000 90.300 97.400 90.700 ;
        RECT 97.700 90.300 98.100 90.700 ;
        RECT 97.000 70.300 97.400 70.700 ;
        RECT 97.700 70.300 98.100 70.700 ;
        RECT 97.000 50.300 97.400 50.700 ;
        RECT 97.700 50.300 98.100 50.700 ;
        RECT 97.000 30.300 97.400 30.700 ;
        RECT 97.700 30.300 98.100 30.700 ;
        RECT 97.000 10.300 97.400 10.700 ;
        RECT 97.700 10.300 98.100 10.700 ;
      LAYER metal3 ;
        RECT 96.800 170.300 98.400 170.700 ;
        RECT 96.800 150.300 98.400 150.700 ;
        RECT 96.800 130.300 98.400 130.700 ;
        RECT 96.800 110.300 98.400 110.700 ;
        RECT 96.800 90.300 98.400 90.700 ;
        RECT 96.800 70.300 98.400 70.700 ;
        RECT 96.800 50.300 98.400 50.700 ;
        RECT 96.800 30.300 98.400 30.700 ;
        RECT 96.800 10.300 98.400 10.700 ;
      LAYER via3 ;
        RECT 97.000 170.300 97.400 170.700 ;
        RECT 97.800 170.300 98.200 170.700 ;
        RECT 97.000 150.300 97.400 150.700 ;
        RECT 97.800 150.300 98.200 150.700 ;
        RECT 97.000 130.300 97.400 130.700 ;
        RECT 97.800 130.300 98.200 130.700 ;
        RECT 97.000 110.300 97.400 110.700 ;
        RECT 97.800 110.300 98.200 110.700 ;
        RECT 97.000 90.300 97.400 90.700 ;
        RECT 97.800 90.300 98.200 90.700 ;
        RECT 97.000 70.300 97.400 70.700 ;
        RECT 97.800 70.300 98.200 70.700 ;
        RECT 97.000 50.300 97.400 50.700 ;
        RECT 97.800 50.300 98.200 50.700 ;
        RECT 97.000 30.300 97.400 30.700 ;
        RECT 97.800 30.300 98.200 30.700 ;
        RECT 97.000 10.300 97.400 10.700 ;
        RECT 97.800 10.300 98.200 10.700 ;
      LAYER metal4 ;
        RECT 96.800 170.300 98.400 170.700 ;
        RECT 96.800 150.300 98.400 150.700 ;
        RECT 96.800 130.300 98.400 130.700 ;
        RECT 96.800 110.300 98.400 110.700 ;
        RECT 96.800 90.300 98.400 90.700 ;
        RECT 96.800 70.300 98.400 70.700 ;
        RECT 96.800 50.300 98.400 50.700 ;
        RECT 96.800 30.300 98.400 30.700 ;
        RECT 96.800 10.300 98.400 10.700 ;
      LAYER via4 ;
        RECT 97.000 170.300 97.400 170.700 ;
        RECT 97.700 170.300 98.100 170.700 ;
        RECT 97.000 150.300 97.400 150.700 ;
        RECT 97.700 150.300 98.100 150.700 ;
        RECT 97.000 130.300 97.400 130.700 ;
        RECT 97.700 130.300 98.100 130.700 ;
        RECT 97.000 110.300 97.400 110.700 ;
        RECT 97.700 110.300 98.100 110.700 ;
        RECT 97.000 90.300 97.400 90.700 ;
        RECT 97.700 90.300 98.100 90.700 ;
        RECT 97.000 70.300 97.400 70.700 ;
        RECT 97.700 70.300 98.100 70.700 ;
        RECT 97.000 50.300 97.400 50.700 ;
        RECT 97.700 50.300 98.100 50.700 ;
        RECT 97.000 30.300 97.400 30.700 ;
        RECT 97.700 30.300 98.100 30.700 ;
        RECT 97.000 10.300 97.400 10.700 ;
        RECT 97.700 10.300 98.100 10.700 ;
      LAYER metal5 ;
        RECT 96.800 170.200 98.400 170.700 ;
        RECT 96.800 150.200 98.400 150.700 ;
        RECT 96.800 130.200 98.400 130.700 ;
        RECT 96.800 110.200 98.400 110.700 ;
        RECT 96.800 90.200 98.400 90.700 ;
        RECT 96.800 70.200 98.400 70.700 ;
        RECT 96.800 50.200 98.400 50.700 ;
        RECT 96.800 30.200 98.400 30.700 ;
        RECT 96.800 10.200 98.400 10.700 ;
      LAYER via5 ;
        RECT 97.800 170.200 98.300 170.700 ;
        RECT 97.800 150.200 98.300 150.700 ;
        RECT 97.800 130.200 98.300 130.700 ;
        RECT 97.800 110.200 98.300 110.700 ;
        RECT 97.800 90.200 98.300 90.700 ;
        RECT 97.800 70.200 98.300 70.700 ;
        RECT 97.800 50.200 98.300 50.700 ;
        RECT 97.800 30.200 98.300 30.700 ;
        RECT 97.800 10.200 98.300 10.700 ;
      LAYER metal6 ;
        RECT 96.800 -3.000 98.400 173.000 ;
    END
  END gnd
  PIN clock
    PORT
      LAYER metal1 ;
        RECT 82.200 106.900 82.600 107.200 ;
        RECT 122.200 106.900 122.600 107.200 ;
        RECT 81.700 106.500 82.600 106.900 ;
        RECT 121.700 106.500 122.600 106.900 ;
        RECT 175.000 106.900 175.400 107.200 ;
        RECT 175.000 106.500 175.900 106.900 ;
        RECT 99.000 94.100 99.900 94.500 ;
        RECT 99.000 93.800 99.400 94.100 ;
        RECT 63.800 46.900 64.200 47.200 ;
        RECT 63.300 46.500 64.200 46.900 ;
        RECT 139.000 34.100 139.900 34.500 ;
        RECT 139.000 33.800 139.400 34.100 ;
        RECT 129.400 26.900 129.800 27.200 ;
        RECT 128.900 26.500 129.800 26.900 ;
        RECT 64.900 14.100 65.800 14.500 ;
        RECT 65.400 13.800 65.800 14.100 ;
      LAYER via1 ;
        RECT 82.200 106.800 82.600 107.200 ;
        RECT 122.200 106.800 122.600 107.200 ;
        RECT 175.000 106.800 175.400 107.200 ;
        RECT 63.800 46.800 64.200 47.200 ;
        RECT 129.400 26.800 129.800 27.200 ;
      LAYER metal2 ;
        RECT 82.200 106.800 82.600 107.200 ;
        RECT 122.200 106.800 122.600 107.200 ;
        RECT 175.000 106.800 175.400 107.200 ;
        RECT 82.200 100.200 82.500 106.800 ;
        RECT 122.200 105.200 122.500 106.800 ;
        RECT 175.000 105.200 175.300 106.800 ;
        RECT 122.200 104.800 122.600 105.200 ;
        RECT 175.000 104.800 175.400 105.200 ;
        RECT 122.200 100.200 122.500 104.800 ;
        RECT 82.200 99.800 82.600 100.200 ;
        RECT 99.000 99.800 99.400 100.200 ;
        RECT 122.200 99.800 122.600 100.200 ;
        RECT 99.000 94.200 99.300 99.800 ;
        RECT 99.000 93.800 99.400 94.200 ;
        RECT 63.800 47.800 64.200 48.200 ;
        RECT 63.800 47.200 64.100 47.800 ;
        RECT 63.800 46.800 64.200 47.200 ;
        RECT 139.000 34.800 139.400 35.200 ;
        RECT 139.000 34.200 139.300 34.800 ;
        RECT 139.000 33.800 139.400 34.200 ;
        RECT 139.000 27.200 139.300 33.800 ;
        RECT 128.600 27.100 129.000 27.200 ;
        RECT 129.400 27.100 129.800 27.200 ;
        RECT 128.600 26.800 129.800 27.100 ;
        RECT 139.000 26.800 139.400 27.200 ;
        RECT 64.600 14.100 65.000 14.200 ;
        RECT 65.400 14.100 65.800 14.200 ;
        RECT 64.600 13.800 65.800 14.100 ;
        RECT 65.400 -1.800 65.700 13.800 ;
        RECT 65.400 -2.200 65.800 -1.800 ;
      LAYER metal3 ;
        RECT 122.200 105.100 122.600 105.200 ;
        RECT 139.000 105.100 139.400 105.200 ;
        RECT 175.000 105.100 175.400 105.200 ;
        RECT 122.200 104.800 175.400 105.100 ;
        RECT 64.600 100.100 65.000 100.200 ;
        RECT 82.200 100.100 82.600 100.200 ;
        RECT 99.000 100.100 99.400 100.200 ;
        RECT 122.200 100.100 122.600 100.200 ;
        RECT 64.600 99.800 122.600 100.100 ;
        RECT 63.800 47.800 64.200 48.200 ;
        RECT 63.800 47.100 64.100 47.800 ;
        RECT 64.600 47.100 65.000 47.200 ;
        RECT 63.800 46.800 65.000 47.100 ;
        RECT 139.000 34.800 139.400 35.200 ;
        RECT 139.000 34.200 139.300 34.800 ;
        RECT 139.000 33.800 139.400 34.200 ;
        RECT 128.600 27.100 129.000 27.200 ;
        RECT 139.000 27.100 139.400 27.200 ;
        RECT 128.600 26.800 139.400 27.100 ;
        RECT 64.600 14.100 65.000 14.200 ;
        RECT 65.400 14.100 65.800 14.200 ;
        RECT 64.600 13.800 65.800 14.100 ;
      LAYER via3 ;
        RECT 139.000 104.800 139.400 105.200 ;
        RECT 64.600 46.800 65.000 47.200 ;
        RECT 65.400 13.800 65.800 14.200 ;
      LAYER metal4 ;
        RECT 139.000 104.800 139.400 105.200 ;
        RECT 64.600 99.800 65.000 100.200 ;
        RECT 64.600 47.200 64.900 99.800 ;
        RECT 64.600 46.800 65.000 47.200 ;
        RECT 64.600 14.100 64.900 46.800 ;
        RECT 139.000 34.200 139.300 104.800 ;
        RECT 139.000 33.800 139.400 34.200 ;
        RECT 65.400 14.100 65.800 14.200 ;
        RECT 64.600 13.800 65.800 14.100 ;
    END
  END clock
  PIN key[0]
    PORT
      LAYER metal1 ;
        RECT 169.400 154.800 169.800 155.600 ;
        RECT 169.400 147.800 169.800 148.600 ;
      LAYER metal2 ;
        RECT 170.200 172.800 170.600 173.200 ;
        RECT 170.200 170.200 170.500 172.800 ;
        RECT 168.600 169.800 169.000 170.200 ;
        RECT 170.200 169.800 170.600 170.200 ;
        RECT 168.600 155.100 168.900 169.800 ;
        RECT 169.400 155.100 169.800 155.200 ;
        RECT 168.600 154.800 169.800 155.100 ;
        RECT 169.400 148.200 169.700 154.800 ;
        RECT 169.400 147.800 169.800 148.200 ;
      LAYER metal3 ;
        RECT 168.600 170.100 169.000 170.200 ;
        RECT 170.200 170.100 170.600 170.200 ;
        RECT 168.600 169.800 170.600 170.100 ;
    END
  END key[0]
  PIN key[1]
    PORT
      LAYER metal1 ;
        RECT 166.200 155.100 166.600 155.200 ;
        RECT 165.400 154.800 166.600 155.100 ;
        RECT 176.600 154.800 177.000 155.600 ;
        RECT 165.400 153.800 165.800 154.800 ;
      LAYER via1 ;
        RECT 166.200 154.800 166.600 155.200 ;
      LAYER metal2 ;
        RECT 175.800 173.100 176.200 173.200 ;
        RECT 175.800 172.800 176.900 173.100 ;
        RECT 176.600 156.200 176.900 172.800 ;
        RECT 166.200 155.800 166.600 156.200 ;
        RECT 176.600 155.800 177.000 156.200 ;
        RECT 166.200 155.200 166.500 155.800 ;
        RECT 176.600 155.200 176.900 155.800 ;
        RECT 166.200 154.800 166.600 155.200 ;
        RECT 176.600 154.800 177.000 155.200 ;
      LAYER metal3 ;
        RECT 166.200 156.100 166.600 156.200 ;
        RECT 176.600 156.100 177.000 156.200 ;
        RECT 166.200 155.800 177.000 156.100 ;
    END
  END key[1]
  PIN key[2]
    PORT
      LAYER metal1 ;
        RECT 166.200 146.100 166.600 146.200 ;
        RECT 167.800 146.100 168.200 146.200 ;
        RECT 166.200 145.800 168.200 146.100 ;
        RECT 166.200 145.400 166.600 145.800 ;
        RECT 167.800 145.400 168.200 145.800 ;
      LAYER via1 ;
        RECT 167.800 145.800 168.200 146.200 ;
      LAYER metal2 ;
        RECT 167.800 172.800 168.200 173.200 ;
        RECT 167.800 146.200 168.100 172.800 ;
        RECT 167.800 145.800 168.200 146.200 ;
    END
  END key[2]
  PIN key[3]
    PORT
      LAYER metal1 ;
        RECT 152.600 165.400 153.000 166.200 ;
        RECT 164.600 154.800 165.000 155.200 ;
        RECT 164.600 154.400 164.900 154.800 ;
        RECT 164.400 154.100 164.900 154.400 ;
        RECT 164.400 154.000 164.800 154.100 ;
      LAYER via1 ;
        RECT 152.600 165.800 153.000 166.200 ;
      LAYER metal2 ;
        RECT 151.000 172.800 151.400 173.200 ;
        RECT 151.000 170.200 151.300 172.800 ;
        RECT 151.000 169.800 151.400 170.200 ;
        RECT 152.600 169.800 153.000 170.200 ;
        RECT 152.600 166.200 152.900 169.800 ;
        RECT 152.600 165.800 153.000 166.200 ;
        RECT 152.600 165.200 152.900 165.800 ;
        RECT 152.600 164.800 153.000 165.200 ;
        RECT 164.600 164.800 165.000 165.200 ;
        RECT 164.600 155.200 164.900 164.800 ;
        RECT 164.600 154.800 165.000 155.200 ;
      LAYER metal3 ;
        RECT 151.000 170.100 151.400 170.200 ;
        RECT 152.600 170.100 153.000 170.200 ;
        RECT 151.000 169.800 153.000 170.100 ;
        RECT 152.600 165.100 153.000 165.200 ;
        RECT 164.600 165.100 165.000 165.200 ;
        RECT 152.600 164.800 165.000 165.100 ;
    END
  END key[3]
  PIN reset
    PORT
      LAYER metal1 ;
        RECT 131.800 146.900 132.200 147.200 ;
        RECT 131.300 146.500 132.200 146.900 ;
        RECT 142.200 146.900 142.600 147.200 ;
        RECT 142.200 146.500 143.100 146.900 ;
        RECT 108.600 126.900 109.000 127.200 ;
        RECT 108.100 126.500 109.000 126.900 ;
        RECT 122.200 126.900 122.600 127.200 ;
        RECT 122.200 126.500 123.100 126.900 ;
        RECT 0.600 74.100 1.500 74.500 ;
        RECT 127.800 74.100 128.700 74.500 ;
        RECT 0.600 73.800 1.000 74.100 ;
        RECT 127.800 73.800 128.200 74.100 ;
        RECT 3.000 66.900 3.400 67.200 ;
        RECT 123.800 66.900 124.200 67.200 ;
        RECT 140.600 66.900 141.000 67.200 ;
        RECT 3.000 66.500 3.900 66.900 ;
        RECT 123.800 66.500 124.700 66.900 ;
        RECT 140.600 66.500 141.500 66.900 ;
        RECT 0.600 54.100 1.500 54.500 ;
        RECT 0.600 53.800 1.000 54.100 ;
      LAYER via1 ;
        RECT 131.800 146.800 132.200 147.200 ;
        RECT 142.200 146.800 142.600 147.200 ;
        RECT 108.600 126.800 109.000 127.200 ;
        RECT 122.200 126.800 122.600 127.200 ;
        RECT 3.000 66.800 3.400 67.200 ;
        RECT 123.800 66.800 124.200 67.200 ;
        RECT 140.600 66.800 141.000 67.200 ;
      LAYER metal2 ;
        RECT 131.800 146.800 132.200 147.200 ;
        RECT 142.200 146.800 142.600 147.200 ;
        RECT 131.800 144.200 132.100 146.800 ;
        RECT 142.200 144.200 142.500 146.800 ;
        RECT 131.800 143.800 132.200 144.200 ;
        RECT 142.200 143.800 142.600 144.200 ;
        RECT 108.600 127.100 109.000 127.200 ;
        RECT 109.400 127.100 109.800 127.200 ;
        RECT 108.600 126.800 109.800 127.100 ;
        RECT 122.200 127.100 122.600 127.200 ;
        RECT 123.000 127.100 123.400 127.200 ;
        RECT 122.200 126.800 123.400 127.100 ;
        RECT 0.600 74.800 1.000 75.200 ;
        RECT 0.600 74.200 0.900 74.800 ;
        RECT 0.600 73.800 1.000 74.200 ;
        RECT 3.000 73.800 3.400 74.200 ;
        RECT 123.800 73.800 124.200 74.200 ;
        RECT 127.800 74.100 128.200 74.200 ;
        RECT 128.600 74.100 129.000 74.200 ;
        RECT 127.800 73.800 129.000 74.100 ;
        RECT 3.000 67.200 3.300 73.800 ;
        RECT 123.800 67.200 124.100 73.800 ;
        RECT 3.000 66.800 3.400 67.200 ;
        RECT 123.800 66.800 124.200 67.200 ;
        RECT 140.600 66.800 141.000 67.200 ;
        RECT 3.000 63.200 3.300 66.800 ;
        RECT 123.800 63.200 124.100 66.800 ;
        RECT 140.600 63.200 140.900 66.800 ;
        RECT 3.000 62.800 3.400 63.200 ;
        RECT 123.800 62.800 124.200 63.200 ;
        RECT 140.600 62.800 141.000 63.200 ;
        RECT 3.000 54.200 3.300 62.800 ;
        RECT 0.600 54.100 1.000 54.200 ;
        RECT 1.400 54.100 1.800 54.200 ;
        RECT 0.600 53.800 1.800 54.100 ;
        RECT 3.000 53.800 3.400 54.200 ;
      LAYER via2 ;
        RECT 109.400 126.800 109.800 127.200 ;
        RECT 123.000 126.800 123.400 127.200 ;
        RECT 128.600 73.800 129.000 74.200 ;
        RECT 1.400 53.800 1.800 54.200 ;
      LAYER metal3 ;
        RECT 122.200 144.100 122.600 144.200 ;
        RECT 131.800 144.100 132.200 144.200 ;
        RECT 142.200 144.100 142.600 144.200 ;
        RECT 122.200 143.800 142.600 144.100 ;
        RECT 109.400 127.100 109.800 127.200 ;
        RECT 122.200 127.100 122.600 127.200 ;
        RECT 123.000 127.100 123.400 127.200 ;
        RECT 109.400 126.800 123.400 127.100 ;
        RECT 0.600 74.800 1.000 75.200 ;
        RECT -2.600 74.100 -2.200 74.200 ;
        RECT 0.600 74.100 0.900 74.800 ;
        RECT 3.000 74.100 3.400 74.200 ;
        RECT -2.600 73.800 3.400 74.100 ;
        RECT 122.200 74.100 122.600 74.200 ;
        RECT 123.800 74.100 124.200 74.200 ;
        RECT 128.600 74.100 129.000 74.200 ;
        RECT 122.200 73.800 129.000 74.100 ;
        RECT 3.000 63.100 3.400 63.200 ;
        RECT 123.800 63.100 124.200 63.200 ;
        RECT 140.600 63.100 141.000 63.200 ;
        RECT 3.000 62.800 141.000 63.100 ;
        RECT 1.400 54.100 1.800 54.200 ;
        RECT 3.000 54.100 3.400 54.200 ;
        RECT 1.400 53.800 3.400 54.100 ;
      LAYER via3 ;
        RECT 122.200 126.800 122.600 127.200 ;
      LAYER metal4 ;
        RECT 122.200 143.800 122.600 144.200 ;
        RECT 122.200 127.200 122.500 143.800 ;
        RECT 122.200 126.800 122.600 127.200 ;
        RECT 122.200 74.200 122.500 126.800 ;
        RECT 122.200 73.800 122.600 74.200 ;
    END
  END reset
  PIN time_button
    PORT
      LAYER metal1 ;
        RECT 0.600 27.800 1.000 28.600 ;
        RECT 7.000 27.800 7.400 28.600 ;
        RECT 3.800 27.100 4.200 27.200 ;
        RECT 4.600 27.100 5.100 27.200 ;
        RECT 3.800 26.800 5.100 27.100 ;
        RECT 4.800 26.400 5.200 26.800 ;
      LAYER metal2 ;
        RECT 0.600 27.800 1.000 28.200 ;
        RECT 7.000 27.800 7.400 28.200 ;
        RECT 0.600 25.200 0.900 27.800 ;
        RECT 3.800 26.800 4.200 27.200 ;
        RECT 3.800 25.200 4.100 26.800 ;
        RECT 7.000 25.200 7.300 27.800 ;
        RECT 0.600 24.800 1.000 25.200 ;
        RECT 3.800 24.800 4.200 25.200 ;
        RECT 7.000 24.800 7.400 25.200 ;
      LAYER metal3 ;
        RECT -2.600 25.100 -2.200 25.200 ;
        RECT 0.600 25.100 1.000 25.200 ;
        RECT 3.800 25.100 4.200 25.200 ;
        RECT 7.000 25.100 7.400 25.200 ;
        RECT -2.600 24.800 7.400 25.100 ;
    END
  END time_button
  PIN alarm_button
    PORT
      LAYER metal1 ;
        RECT 65.400 32.400 65.800 33.200 ;
        RECT 67.800 32.400 68.200 33.200 ;
        RECT 75.800 32.400 76.200 33.200 ;
        RECT 68.600 27.800 69.000 28.600 ;
        RECT 76.600 26.800 77.000 27.600 ;
      LAYER via1 ;
        RECT 65.400 32.800 65.800 33.200 ;
        RECT 67.800 32.800 68.200 33.200 ;
        RECT 75.800 32.800 76.200 33.200 ;
      LAYER metal2 ;
        RECT 65.400 32.800 65.800 33.200 ;
        RECT 67.800 32.800 68.200 33.200 ;
        RECT 75.800 32.800 76.200 33.200 ;
        RECT 65.400 32.200 65.700 32.800 ;
        RECT 65.400 31.800 65.800 32.200 ;
        RECT 67.800 29.100 68.100 32.800 ;
        RECT 75.800 31.100 76.100 32.800 ;
        RECT 75.800 30.800 76.900 31.100 ;
        RECT 68.600 29.100 69.000 29.200 ;
        RECT 67.800 28.800 69.000 29.100 ;
        RECT 68.600 28.200 68.900 28.800 ;
        RECT 76.600 28.200 76.900 30.800 ;
        RECT 68.600 27.800 69.000 28.200 ;
        RECT 76.600 27.800 77.000 28.200 ;
        RECT 76.600 27.200 76.900 27.800 ;
        RECT 76.600 26.800 77.000 27.200 ;
        RECT 76.600 1.800 77.000 2.200 ;
        RECT 76.600 -1.800 76.900 1.800 ;
        RECT 76.600 -2.200 77.000 -1.800 ;
      LAYER via2 ;
        RECT 68.600 28.800 69.000 29.200 ;
      LAYER metal3 ;
        RECT 67.800 33.100 68.200 33.200 ;
        RECT 65.400 32.800 68.200 33.100 ;
        RECT 65.400 32.200 65.700 32.800 ;
        RECT 65.400 31.800 65.800 32.200 ;
        RECT 68.600 28.800 69.000 29.200 ;
        RECT 68.600 28.100 68.900 28.800 ;
        RECT 76.600 28.100 77.000 28.200 ;
        RECT 68.600 27.800 77.000 28.100 ;
        RECT 76.600 2.800 77.000 3.200 ;
        RECT 76.600 2.200 76.900 2.800 ;
        RECT 76.600 1.800 77.000 2.200 ;
      LAYER via3 ;
        RECT 76.600 27.800 77.000 28.200 ;
      LAYER metal4 ;
        RECT 76.600 27.800 77.000 28.200 ;
        RECT 76.600 3.200 76.900 27.800 ;
        RECT 76.600 2.800 77.000 3.200 ;
    END
  END alarm_button
  PIN fastwatch
    PORT
      LAYER metal1 ;
        RECT 158.200 85.800 158.600 86.600 ;
        RECT 160.600 84.400 161.000 85.200 ;
      LAYER via1 ;
        RECT 160.600 84.800 161.000 85.200 ;
      LAYER metal2 ;
        RECT 158.200 86.100 158.600 86.200 ;
        RECT 159.000 86.100 159.400 86.200 ;
        RECT 158.200 85.800 159.400 86.100 ;
        RECT 160.600 85.800 161.000 86.200 ;
        RECT 160.600 85.200 160.900 85.800 ;
        RECT 160.600 84.800 161.000 85.200 ;
      LAYER via2 ;
        RECT 159.000 85.800 159.400 86.200 ;
      LAYER metal3 ;
        RECT 159.000 86.100 159.400 86.200 ;
        RECT 160.600 86.100 161.000 86.200 ;
        RECT 164.600 86.100 165.000 86.200 ;
        RECT 159.000 85.800 165.000 86.100 ;
        RECT 186.200 85.100 186.600 85.200 ;
        RECT 198.200 85.100 198.600 85.200 ;
        RECT 186.200 84.800 198.600 85.100 ;
      LAYER via3 ;
        RECT 164.600 85.800 165.000 86.200 ;
      LAYER metal4 ;
        RECT 164.600 85.800 165.000 86.200 ;
        RECT 164.600 85.200 164.900 85.800 ;
        RECT 164.600 84.800 165.000 85.200 ;
        RECT 185.400 85.100 185.800 85.200 ;
        RECT 186.200 85.100 186.600 85.200 ;
        RECT 185.400 84.800 186.600 85.100 ;
      LAYER metal5 ;
        RECT 164.600 85.100 165.000 85.200 ;
        RECT 185.400 85.100 185.800 85.200 ;
        RECT 164.600 84.800 185.800 85.100 ;
    END
  END fastwatch
  PIN ms_hour[0]
    PORT
      LAYER metal1 ;
        RECT 22.200 166.200 22.600 169.900 ;
        RECT 22.300 165.100 22.600 166.200 ;
        RECT 22.200 161.100 22.600 165.100 ;
      LAYER via1 ;
        RECT 22.200 168.800 22.600 169.200 ;
      LAYER metal2 ;
        RECT 21.400 173.100 21.800 173.200 ;
        RECT 21.400 172.800 22.500 173.100 ;
        RECT 22.200 169.200 22.500 172.800 ;
        RECT 22.200 168.800 22.600 169.200 ;
    END
  END ms_hour[0]
  PIN ms_hour[1]
    PORT
      LAYER metal1 ;
        RECT 17.400 166.200 17.800 169.900 ;
        RECT 17.500 165.100 17.800 166.200 ;
        RECT 17.400 161.100 17.800 165.100 ;
      LAYER via1 ;
        RECT 17.400 168.800 17.800 169.200 ;
      LAYER metal2 ;
        RECT 16.600 173.100 17.000 173.200 ;
        RECT 16.600 172.800 17.700 173.100 ;
        RECT 17.400 169.200 17.700 172.800 ;
        RECT 17.400 168.800 17.800 169.200 ;
    END
  END ms_hour[1]
  PIN ms_hour[2]
    PORT
      LAYER metal1 ;
        RECT 0.600 166.200 1.000 169.900 ;
        RECT 0.600 165.100 0.900 166.200 ;
        RECT 0.600 161.100 1.000 165.100 ;
      LAYER via1 ;
        RECT 0.600 166.800 1.000 167.200 ;
      LAYER metal2 ;
        RECT 0.600 167.800 1.000 168.200 ;
        RECT 0.600 167.200 0.900 167.800 ;
        RECT 0.600 166.800 1.000 167.200 ;
      LAYER metal3 ;
        RECT 0.600 167.800 1.000 168.200 ;
        RECT -2.600 167.100 -2.200 167.200 ;
        RECT 0.600 167.100 0.900 167.800 ;
        RECT -2.600 166.800 0.900 167.100 ;
    END
  END ms_hour[2]
  PIN ms_hour[3]
    PORT
      LAYER metal1 ;
        RECT 3.000 166.200 3.400 169.900 ;
        RECT 3.000 165.100 3.300 166.200 ;
        RECT 3.000 161.100 3.400 165.100 ;
      LAYER via1 ;
        RECT 3.000 166.800 3.400 167.200 ;
      LAYER metal2 ;
        RECT 3.000 166.800 3.400 167.200 ;
        RECT 3.000 165.200 3.300 166.800 ;
        RECT 3.000 164.800 3.400 165.200 ;
      LAYER metal3 ;
        RECT -2.600 165.100 -2.200 165.200 ;
        RECT 3.000 165.100 3.400 165.200 ;
        RECT -2.600 164.800 3.400 165.100 ;
    END
  END ms_hour[3]
  PIN ms_hour[4]
    PORT
      LAYER metal1 ;
        RECT 175.000 166.200 175.400 169.900 ;
        RECT 175.100 165.100 175.400 166.200 ;
        RECT 175.000 161.100 175.400 165.100 ;
      LAYER via1 ;
        RECT 175.000 168.800 175.400 169.200 ;
      LAYER metal2 ;
        RECT 174.200 173.100 174.600 173.200 ;
        RECT 174.200 172.800 175.300 173.100 ;
        RECT 175.000 169.200 175.300 172.800 ;
        RECT 175.000 168.800 175.400 169.200 ;
    END
  END ms_hour[4]
  PIN ms_hour[5]
    PORT
      LAYER metal1 ;
        RECT 191.000 66.200 191.400 69.900 ;
        RECT 191.100 65.100 191.400 66.200 ;
        RECT 191.000 61.100 191.400 65.100 ;
      LAYER via1 ;
        RECT 191.000 63.800 191.400 64.200 ;
      LAYER metal2 ;
        RECT 191.000 64.800 191.400 65.200 ;
        RECT 191.000 64.200 191.300 64.800 ;
        RECT 191.000 63.800 191.400 64.200 ;
      LAYER metal3 ;
        RECT 191.000 65.100 191.400 65.200 ;
        RECT 198.200 65.100 198.600 65.200 ;
        RECT 191.000 64.800 198.600 65.100 ;
    END
  END ms_hour[5]
  PIN ms_hour[6]
    PORT
      LAYER metal1 ;
        RECT 0.600 66.200 1.000 69.900 ;
        RECT 0.600 65.100 0.900 66.200 ;
        RECT 0.600 61.100 1.000 65.100 ;
      LAYER via1 ;
        RECT 0.600 63.800 1.000 64.200 ;
      LAYER metal2 ;
        RECT 0.600 64.800 1.000 65.200 ;
        RECT 0.600 64.200 0.900 64.800 ;
        RECT 0.600 63.800 1.000 64.200 ;
      LAYER metal3 ;
        RECT -2.600 65.100 -2.200 65.200 ;
        RECT 0.600 65.100 1.000 65.200 ;
        RECT -2.600 64.800 1.000 65.100 ;
    END
  END ms_hour[6]
  PIN ms_hour[7]
    PORT
      LAYER metal1 ;
        RECT 0.600 46.200 1.000 49.900 ;
        RECT 0.600 45.100 0.900 46.200 ;
        RECT 0.600 41.100 1.000 45.100 ;
      LAYER via1 ;
        RECT 0.600 43.800 1.000 44.200 ;
      LAYER metal2 ;
        RECT 0.600 44.800 1.000 45.200 ;
        RECT 0.600 44.200 0.900 44.800 ;
        RECT 0.600 43.800 1.000 44.200 ;
      LAYER metal3 ;
        RECT -2.600 45.100 -2.200 45.200 ;
        RECT 0.600 45.100 1.000 45.200 ;
        RECT -2.600 44.800 1.000 45.100 ;
    END
  END ms_hour[7]
  PIN ls_hour[0]
    PORT
      LAYER metal1 ;
        RECT 107.000 155.900 107.400 159.900 ;
        RECT 107.100 154.800 107.400 155.900 ;
        RECT 107.000 151.100 107.400 154.800 ;
      LAYER via1 ;
        RECT 107.000 158.800 107.400 159.200 ;
      LAYER metal2 ;
        RECT 106.200 172.800 106.600 173.200 ;
        RECT 106.200 170.200 106.500 172.800 ;
        RECT 106.200 169.800 106.600 170.200 ;
        RECT 107.000 160.800 107.400 161.200 ;
        RECT 107.000 159.200 107.300 160.800 ;
        RECT 107.000 158.800 107.400 159.200 ;
      LAYER metal3 ;
        RECT 106.200 170.100 106.600 170.200 ;
        RECT 107.000 170.100 107.400 170.200 ;
        RECT 106.200 169.800 107.400 170.100 ;
        RECT 106.200 161.100 106.600 161.200 ;
        RECT 107.000 161.100 107.400 161.200 ;
        RECT 106.200 160.800 107.400 161.100 ;
      LAYER via3 ;
        RECT 107.000 169.800 107.400 170.200 ;
      LAYER metal4 ;
        RECT 107.000 170.100 107.400 170.200 ;
        RECT 106.200 169.800 107.400 170.100 ;
        RECT 106.200 161.200 106.500 169.800 ;
        RECT 106.200 160.800 106.600 161.200 ;
    END
  END ls_hour[0]
  PIN ls_hour[1]
    PORT
      LAYER metal1 ;
        RECT 109.400 155.900 109.800 159.900 ;
        RECT 109.500 154.800 109.800 155.900 ;
        RECT 109.400 151.100 109.800 154.800 ;
      LAYER via1 ;
        RECT 109.400 158.800 109.800 159.200 ;
      LAYER metal2 ;
        RECT 109.400 173.100 109.800 173.200 ;
        RECT 109.400 172.800 110.500 173.100 ;
        RECT 110.200 162.100 110.500 172.800 ;
        RECT 109.400 161.800 110.500 162.100 ;
        RECT 109.400 159.200 109.700 161.800 ;
        RECT 109.400 158.800 109.800 159.200 ;
    END
  END ls_hour[1]
  PIN ls_hour[2]
    PORT
      LAYER metal1 ;
        RECT 82.200 166.200 82.600 169.900 ;
        RECT 82.200 165.100 82.500 166.200 ;
        RECT 82.200 161.100 82.600 165.100 ;
      LAYER via1 ;
        RECT 82.200 168.800 82.600 169.200 ;
      LAYER metal2 ;
        RECT 83.000 173.100 83.400 173.200 ;
        RECT 82.200 172.800 83.400 173.100 ;
        RECT 82.200 169.200 82.500 172.800 ;
        RECT 82.200 168.800 82.600 169.200 ;
    END
  END ls_hour[2]
  PIN ls_hour[3]
    PORT
      LAYER metal1 ;
        RECT 87.000 166.200 87.400 169.900 ;
        RECT 87.000 165.100 87.300 166.200 ;
        RECT 87.000 161.100 87.400 165.100 ;
      LAYER via1 ;
        RECT 87.000 168.800 87.400 169.200 ;
      LAYER metal2 ;
        RECT 87.800 173.100 88.200 173.200 ;
        RECT 87.000 172.800 88.200 173.100 ;
        RECT 87.000 169.200 87.300 172.800 ;
        RECT 87.000 168.800 87.400 169.200 ;
    END
  END ls_hour[3]
  PIN ls_hour[4]
    PORT
      LAYER metal1 ;
        RECT 131.000 166.200 131.400 169.900 ;
        RECT 131.000 165.100 131.300 166.200 ;
        RECT 131.000 161.100 131.400 165.100 ;
      LAYER via1 ;
        RECT 131.000 168.800 131.400 169.200 ;
      LAYER metal2 ;
        RECT 131.000 172.800 131.400 173.200 ;
        RECT 131.000 169.200 131.300 172.800 ;
        RECT 131.000 168.800 131.400 169.200 ;
    END
  END ls_hour[4]
  PIN ls_hour[5]
    PORT
      LAYER metal1 ;
        RECT 191.800 166.200 192.200 169.900 ;
        RECT 191.900 165.100 192.200 166.200 ;
        RECT 191.800 161.100 192.200 165.100 ;
      LAYER via1 ;
        RECT 191.800 168.800 192.200 169.200 ;
      LAYER metal2 ;
        RECT 191.000 173.100 191.400 173.200 ;
        RECT 191.000 172.800 192.100 173.100 ;
        RECT 191.800 169.200 192.100 172.800 ;
        RECT 191.800 168.800 192.200 169.200 ;
    END
  END ls_hour[5]
  PIN ls_hour[6]
    PORT
      LAYER metal1 ;
        RECT 106.200 166.200 106.600 169.900 ;
        RECT 106.300 165.100 106.600 166.200 ;
        RECT 106.200 161.100 106.600 165.100 ;
      LAYER via1 ;
        RECT 106.200 168.800 106.600 169.200 ;
      LAYER metal2 ;
        RECT 107.800 172.800 108.200 173.200 ;
        RECT 107.800 169.200 108.100 172.800 ;
        RECT 106.200 168.800 106.600 169.200 ;
        RECT 107.800 168.800 108.200 169.200 ;
        RECT 106.200 168.200 106.500 168.800 ;
        RECT 106.200 167.800 106.600 168.200 ;
      LAYER metal3 ;
        RECT 107.800 169.100 108.200 169.200 ;
        RECT 106.200 168.800 108.200 169.100 ;
        RECT 106.200 168.200 106.500 168.800 ;
        RECT 106.200 167.800 106.600 168.200 ;
    END
  END ls_hour[6]
  PIN ls_hour[7]
    PORT
      LAYER metal1 ;
        RECT 191.000 135.900 191.400 139.900 ;
        RECT 191.100 134.800 191.400 135.900 ;
        RECT 191.000 131.100 191.400 134.800 ;
      LAYER via1 ;
        RECT 191.000 136.800 191.400 137.200 ;
      LAYER metal2 ;
        RECT 191.000 137.800 191.400 138.200 ;
        RECT 191.000 137.200 191.300 137.800 ;
        RECT 191.000 136.800 191.400 137.200 ;
      LAYER metal3 ;
        RECT 191.000 137.800 191.400 138.200 ;
        RECT 191.000 137.100 191.300 137.800 ;
        RECT 198.200 137.100 198.600 137.200 ;
        RECT 191.000 136.800 198.600 137.100 ;
    END
  END ls_hour[7]
  PIN ms_minute[0]
    PORT
      LAYER metal1 ;
        RECT 115.000 155.900 115.400 159.900 ;
        RECT 115.000 154.800 115.300 155.900 ;
        RECT 115.000 151.100 115.400 154.800 ;
      LAYER via1 ;
        RECT 115.000 158.800 115.400 159.200 ;
      LAYER metal2 ;
        RECT 115.800 172.800 116.200 173.200 ;
        RECT 115.800 170.200 116.100 172.800 ;
        RECT 115.800 169.800 116.200 170.200 ;
        RECT 115.000 165.800 115.400 166.200 ;
        RECT 115.000 159.200 115.300 165.800 ;
        RECT 115.000 158.800 115.400 159.200 ;
      LAYER metal3 ;
        RECT 115.000 170.100 115.400 170.200 ;
        RECT 115.800 170.100 116.200 170.200 ;
        RECT 115.000 169.800 116.200 170.100 ;
        RECT 115.000 166.100 115.400 166.200 ;
        RECT 115.800 166.100 116.200 166.200 ;
        RECT 115.000 165.800 116.200 166.100 ;
      LAYER via3 ;
        RECT 115.800 165.800 116.200 166.200 ;
      LAYER metal4 ;
        RECT 115.000 170.100 115.400 170.200 ;
        RECT 115.000 169.800 116.100 170.100 ;
        RECT 115.800 166.200 116.100 169.800 ;
        RECT 115.800 165.800 116.200 166.200 ;
    END
  END ms_minute[0]
  PIN ms_minute[1]
    PORT
      LAYER metal1 ;
        RECT 116.600 166.200 117.000 169.900 ;
        RECT 116.600 165.100 116.900 166.200 ;
        RECT 116.600 161.100 117.000 165.100 ;
      LAYER via1 ;
        RECT 116.600 168.800 117.000 169.200 ;
      LAYER metal2 ;
        RECT 117.400 173.100 117.800 173.200 ;
        RECT 116.600 172.800 117.800 173.100 ;
        RECT 116.600 169.200 116.900 172.800 ;
        RECT 116.600 168.800 117.000 169.200 ;
    END
  END ms_minute[1]
  PIN ms_minute[2]
    PORT
      LAYER metal1 ;
        RECT 131.800 155.900 132.200 159.900 ;
        RECT 131.900 154.800 132.200 155.900 ;
        RECT 131.800 151.100 132.200 154.800 ;
      LAYER via1 ;
        RECT 131.800 158.800 132.200 159.200 ;
      LAYER metal2 ;
        RECT 132.600 172.800 133.000 173.200 ;
        RECT 132.600 170.200 132.900 172.800 ;
        RECT 132.600 169.800 133.000 170.200 ;
        RECT 131.800 162.800 132.200 163.200 ;
        RECT 131.800 159.200 132.100 162.800 ;
        RECT 131.800 158.800 132.200 159.200 ;
      LAYER metal3 ;
        RECT 131.800 170.100 132.200 170.200 ;
        RECT 132.600 170.100 133.000 170.200 ;
        RECT 131.800 169.800 133.000 170.100 ;
        RECT 131.800 163.100 132.200 163.200 ;
        RECT 132.600 163.100 133.000 163.200 ;
        RECT 131.800 162.800 133.000 163.100 ;
      LAYER via3 ;
        RECT 132.600 162.800 133.000 163.200 ;
      LAYER metal4 ;
        RECT 131.800 170.100 132.200 170.200 ;
        RECT 131.800 169.800 132.900 170.100 ;
        RECT 132.600 163.200 132.900 169.800 ;
        RECT 132.600 162.800 133.000 163.200 ;
    END
  END ms_minute[2]
  PIN ms_minute[3]
    PORT
      LAYER metal1 ;
        RECT 120.600 166.200 121.000 169.900 ;
        RECT 120.700 165.100 121.000 166.200 ;
        RECT 120.600 161.100 121.000 165.100 ;
      LAYER via1 ;
        RECT 120.600 168.800 121.000 169.200 ;
      LAYER metal2 ;
        RECT 119.800 173.100 120.200 173.200 ;
        RECT 119.800 172.800 120.900 173.100 ;
        RECT 120.600 169.200 120.900 172.800 ;
        RECT 120.600 168.800 121.000 169.200 ;
    END
  END ms_minute[3]
  PIN ms_minute[4]
    PORT
      LAYER metal1 ;
        RECT 193.400 67.100 193.800 69.900 ;
        RECT 194.200 67.100 194.600 67.200 ;
        RECT 193.400 66.800 194.600 67.100 ;
        RECT 193.400 66.200 193.800 66.800 ;
        RECT 193.500 65.100 193.800 66.200 ;
        RECT 193.400 61.100 193.800 65.100 ;
      LAYER via1 ;
        RECT 194.200 66.800 194.600 67.200 ;
      LAYER metal2 ;
        RECT 194.200 67.100 194.600 67.200 ;
        RECT 195.000 67.100 195.400 67.200 ;
        RECT 194.200 66.800 195.400 67.100 ;
      LAYER via2 ;
        RECT 195.000 66.800 195.400 67.200 ;
      LAYER metal3 ;
        RECT 195.000 67.100 195.400 67.200 ;
        RECT 198.200 67.100 198.600 67.200 ;
        RECT 195.000 66.800 198.600 67.100 ;
    END
  END ms_minute[4]
  PIN ms_minute[5]
    PORT
      LAYER metal1 ;
        RECT 194.200 155.900 194.600 159.900 ;
        RECT 194.300 154.800 194.600 155.900 ;
        RECT 194.200 154.100 194.600 154.800 ;
        RECT 195.000 154.100 195.400 154.200 ;
        RECT 194.200 153.800 195.400 154.100 ;
        RECT 194.200 151.100 194.600 153.800 ;
      LAYER via1 ;
        RECT 195.000 153.800 195.400 154.200 ;
      LAYER metal2 ;
        RECT 195.000 154.800 195.400 155.200 ;
        RECT 195.000 154.200 195.300 154.800 ;
        RECT 195.000 153.800 195.400 154.200 ;
      LAYER metal3 ;
        RECT 195.000 155.100 195.400 155.200 ;
        RECT 198.200 155.100 198.600 155.200 ;
        RECT 195.000 154.800 198.600 155.100 ;
    END
  END ms_minute[5]
  PIN ms_minute[6]
    PORT
      LAYER metal1 ;
        RECT 58.200 6.200 58.600 9.900 ;
        RECT 58.300 5.100 58.600 6.200 ;
        RECT 58.200 1.100 58.600 5.100 ;
      LAYER via1 ;
        RECT 58.200 1.800 58.600 2.200 ;
      LAYER metal2 ;
        RECT 58.200 1.800 58.600 2.200 ;
        RECT 57.400 -1.900 57.800 -1.800 ;
        RECT 58.200 -1.900 58.500 1.800 ;
        RECT 57.400 -2.200 58.500 -1.900 ;
    END
  END ms_minute[6]
  PIN ms_minute[7]
    PORT
      LAYER metal1 ;
        RECT 194.200 95.900 194.600 99.900 ;
        RECT 194.300 94.800 194.600 95.900 ;
        RECT 194.200 91.100 194.600 94.800 ;
      LAYER via1 ;
        RECT 194.200 93.800 194.600 94.200 ;
      LAYER metal2 ;
        RECT 194.200 94.800 194.600 95.200 ;
        RECT 194.200 94.200 194.500 94.800 ;
        RECT 194.200 93.800 194.600 94.200 ;
      LAYER metal3 ;
        RECT 194.200 95.100 194.600 95.200 ;
        RECT 198.200 95.100 198.600 95.200 ;
        RECT 194.200 94.800 198.600 95.100 ;
    END
  END ms_minute[7]
  PIN ls_minute[0]
    PORT
      LAYER metal1 ;
        RECT 192.600 126.200 193.000 129.900 ;
        RECT 192.700 125.100 193.000 126.200 ;
        RECT 192.600 121.100 193.000 125.100 ;
      LAYER via1 ;
        RECT 192.600 123.800 193.000 124.200 ;
      LAYER metal2 ;
        RECT 192.600 124.800 193.000 125.200 ;
        RECT 192.600 124.200 192.900 124.800 ;
        RECT 192.600 123.800 193.000 124.200 ;
      LAYER metal3 ;
        RECT 192.600 125.100 193.000 125.200 ;
        RECT 198.200 125.100 198.600 125.200 ;
        RECT 192.600 124.800 198.600 125.100 ;
    END
  END ls_minute[0]
  PIN ls_minute[1]
    PORT
      LAYER metal1 ;
        RECT 187.800 115.900 188.200 119.900 ;
        RECT 187.900 114.800 188.200 115.900 ;
        RECT 187.800 111.100 188.200 114.800 ;
      LAYER via1 ;
        RECT 187.800 116.800 188.200 117.200 ;
      LAYER metal2 ;
        RECT 187.800 116.800 188.200 117.200 ;
        RECT 187.800 116.200 188.100 116.800 ;
        RECT 187.800 115.800 188.200 116.200 ;
      LAYER metal3 ;
        RECT 187.800 116.100 188.200 116.200 ;
        RECT 187.800 115.800 198.500 116.100 ;
        RECT 198.200 115.200 198.500 115.800 ;
        RECT 198.200 114.800 198.600 115.200 ;
    END
  END ls_minute[1]
  PIN ls_minute[2]
    PORT
      LAYER metal1 ;
        RECT 193.400 87.100 193.800 89.900 ;
        RECT 194.200 87.100 194.600 87.200 ;
        RECT 193.400 86.800 194.600 87.100 ;
        RECT 193.400 86.200 193.800 86.800 ;
        RECT 193.500 85.100 193.800 86.200 ;
        RECT 193.400 81.100 193.800 85.100 ;
      LAYER via1 ;
        RECT 194.200 86.800 194.600 87.200 ;
      LAYER metal2 ;
        RECT 194.200 87.100 194.600 87.200 ;
        RECT 195.000 87.100 195.400 87.200 ;
        RECT 194.200 86.800 195.400 87.100 ;
      LAYER via2 ;
        RECT 195.000 86.800 195.400 87.200 ;
      LAYER metal3 ;
        RECT 195.000 87.100 195.400 87.200 ;
        RECT 198.200 87.100 198.600 87.200 ;
        RECT 195.000 86.800 198.600 87.100 ;
    END
  END ls_minute[2]
  PIN ls_minute[3]
    PORT
      LAYER metal1 ;
        RECT 193.400 135.900 193.800 139.900 ;
        RECT 193.500 134.800 193.800 135.900 ;
        RECT 193.400 134.100 193.800 134.800 ;
        RECT 195.000 134.100 195.400 134.200 ;
        RECT 193.400 133.800 195.400 134.100 ;
        RECT 193.400 131.100 193.800 133.800 ;
      LAYER via1 ;
        RECT 195.000 133.800 195.400 134.200 ;
      LAYER metal2 ;
        RECT 195.000 134.800 195.400 135.200 ;
        RECT 195.000 134.200 195.300 134.800 ;
        RECT 195.000 133.800 195.400 134.200 ;
      LAYER metal3 ;
        RECT 195.000 135.100 195.400 135.200 ;
        RECT 198.200 135.100 198.600 135.200 ;
        RECT 195.000 134.800 198.600 135.100 ;
    END
  END ls_minute[3]
  PIN ls_minute[4]
    PORT
      LAYER metal1 ;
        RECT 189.400 166.200 189.800 169.900 ;
        RECT 189.500 165.100 189.800 166.200 ;
        RECT 189.400 161.100 189.800 165.100 ;
      LAYER via1 ;
        RECT 189.400 168.800 189.800 169.200 ;
      LAYER metal2 ;
        RECT 188.600 173.100 189.000 173.200 ;
        RECT 188.600 172.800 189.700 173.100 ;
        RECT 189.400 169.200 189.700 172.800 ;
        RECT 189.400 168.800 189.800 169.200 ;
    END
  END ls_minute[4]
  PIN ls_minute[5]
    PORT
      LAYER metal1 ;
        RECT 135.000 166.200 135.400 169.900 ;
        RECT 135.100 165.100 135.400 166.200 ;
        RECT 135.000 161.100 135.400 165.100 ;
      LAYER via1 ;
        RECT 135.000 168.800 135.400 169.200 ;
      LAYER metal2 ;
        RECT 134.200 173.100 134.600 173.200 ;
        RECT 134.200 172.800 135.300 173.100 ;
        RECT 135.000 169.200 135.300 172.800 ;
        RECT 135.000 168.800 135.400 169.200 ;
    END
  END ls_minute[5]
  PIN ls_minute[6]
    PORT
      LAYER metal1 ;
        RECT 185.400 166.200 185.800 169.900 ;
        RECT 185.400 165.100 185.700 166.200 ;
        RECT 185.400 161.100 185.800 165.100 ;
      LAYER via1 ;
        RECT 185.400 168.800 185.800 169.200 ;
      LAYER metal2 ;
        RECT 186.200 173.100 186.600 173.200 ;
        RECT 185.400 172.800 186.600 173.100 ;
        RECT 185.400 169.200 185.700 172.800 ;
        RECT 185.400 168.800 185.800 169.200 ;
    END
  END ls_minute[6]
  PIN ls_minute[7]
    PORT
      LAYER metal1 ;
        RECT 0.600 15.900 1.000 19.900 ;
        RECT 0.600 14.800 0.900 15.900 ;
        RECT 0.600 11.100 1.000 14.800 ;
      LAYER via1 ;
        RECT 0.600 13.800 1.000 14.200 ;
      LAYER metal2 ;
        RECT 0.600 14.800 1.000 15.200 ;
        RECT 0.600 14.200 0.900 14.800 ;
        RECT 0.600 13.800 1.000 14.200 ;
      LAYER metal3 ;
        RECT -2.600 15.100 -2.200 15.200 ;
        RECT 0.600 15.100 1.000 15.200 ;
        RECT -2.600 14.800 1.000 15.100 ;
    END
  END ls_minute[7]
  PIN alarm_sound
    PORT
      LAYER metal1 ;
        RECT 0.600 95.900 1.000 99.900 ;
        RECT 0.600 94.800 0.900 95.900 ;
        RECT 0.600 91.100 1.000 94.800 ;
      LAYER via1 ;
        RECT 0.600 93.800 1.000 94.200 ;
      LAYER metal2 ;
        RECT 0.600 94.800 1.000 95.200 ;
        RECT 0.600 94.200 0.900 94.800 ;
        RECT 0.600 93.800 1.000 94.200 ;
      LAYER metal3 ;
        RECT -2.600 95.100 -2.200 95.200 ;
        RECT 0.600 95.100 1.000 95.200 ;
        RECT -2.600 94.800 1.000 95.100 ;
    END
  END alarm_sound
  OBS
      LAYER metal1 ;
        RECT 2.200 167.600 2.600 169.900 ;
        RECT 4.600 167.600 5.000 169.900 ;
        RECT 1.500 167.300 2.600 167.600 ;
        RECT 3.900 167.300 5.000 167.600 ;
        RECT 6.200 168.900 6.600 169.900 ;
        RECT 1.500 165.800 1.800 167.300 ;
        RECT 2.200 165.800 2.600 166.600 ;
        RECT 3.900 165.800 4.200 167.300 ;
        RECT 6.200 167.200 6.500 168.900 ;
        RECT 7.000 167.800 7.400 168.600 ;
        RECT 5.400 166.800 5.800 167.200 ;
        RECT 6.200 166.800 6.600 167.200 ;
        RECT 4.600 166.100 5.000 166.600 ;
        RECT 5.400 166.200 5.700 166.800 ;
        RECT 5.400 166.100 5.800 166.200 ;
        RECT 4.600 165.800 5.800 166.100 ;
        RECT 1.200 165.400 1.800 165.800 ;
        RECT 3.600 165.400 4.200 165.800 ;
        RECT 5.400 165.400 5.800 165.800 ;
        RECT 1.500 165.100 1.800 165.400 ;
        RECT 3.900 165.100 4.200 165.400 ;
        RECT 6.200 165.100 6.500 166.800 ;
        RECT 1.500 164.800 2.600 165.100 ;
        RECT 3.900 164.800 5.000 165.100 ;
        RECT 2.200 161.100 2.600 164.800 ;
        RECT 4.600 161.100 5.000 164.800 ;
        RECT 5.700 164.700 6.600 165.100 ;
        RECT 5.700 161.100 6.100 164.700 ;
        RECT 7.800 161.100 8.200 169.900 ;
        RECT 8.600 167.800 9.000 168.600 ;
        RECT 9.400 168.000 9.800 169.900 ;
        RECT 11.000 168.000 11.400 169.900 ;
        RECT 9.400 167.900 11.400 168.000 ;
        RECT 11.800 167.900 12.200 169.900 ;
        RECT 12.700 168.200 13.100 168.600 ;
        RECT 8.600 167.100 8.900 167.800 ;
        RECT 9.500 167.700 11.300 167.900 ;
        RECT 9.800 167.200 10.200 167.400 ;
        RECT 11.800 167.200 12.100 167.900 ;
        RECT 12.600 167.800 13.000 168.200 ;
        RECT 13.400 167.900 13.800 169.900 ;
        RECT 13.500 167.200 13.800 167.900 ;
        RECT 15.800 167.600 16.200 169.900 ;
        RECT 19.000 168.900 19.400 169.900 ;
        RECT 15.800 167.300 16.900 167.600 ;
        RECT 9.400 167.100 10.200 167.200 ;
        RECT 8.600 166.900 10.200 167.100 ;
        RECT 8.600 166.800 9.800 166.900 ;
        RECT 10.900 166.800 12.200 167.200 ;
        RECT 13.400 166.800 13.800 167.200 ;
        RECT 10.200 165.800 10.600 166.600 ;
        RECT 10.900 165.100 11.200 166.800 ;
        RECT 12.600 166.100 13.000 166.200 ;
        RECT 13.500 166.100 13.800 166.800 ;
        RECT 14.200 166.400 14.600 167.200 ;
        RECT 15.000 166.100 15.400 166.200 ;
        RECT 12.600 165.800 13.800 166.100 ;
        RECT 14.600 165.800 15.400 166.100 ;
        RECT 15.800 165.800 16.200 166.600 ;
        RECT 16.600 165.800 16.900 167.300 ;
        RECT 19.000 167.200 19.300 168.900 ;
        RECT 19.800 167.800 20.200 168.600 ;
        RECT 20.600 167.600 21.000 169.900 ;
        RECT 23.000 167.700 23.400 169.900 ;
        RECT 25.100 169.200 25.700 169.900 ;
        RECT 25.100 168.900 25.800 169.200 ;
        RECT 27.400 168.900 27.800 169.900 ;
        RECT 29.600 169.200 30.000 169.900 ;
        RECT 29.600 168.900 30.600 169.200 ;
        RECT 25.400 168.500 25.800 168.900 ;
        RECT 27.500 168.600 27.800 168.900 ;
        RECT 27.500 168.300 28.900 168.600 ;
        RECT 28.500 168.200 28.900 168.300 ;
        RECT 29.400 168.200 29.800 168.600 ;
        RECT 30.200 168.500 30.600 168.900 ;
        RECT 24.500 167.700 24.900 167.800 ;
        RECT 20.600 167.300 21.700 167.600 ;
        RECT 19.000 166.800 19.400 167.200 ;
        RECT 11.800 165.100 12.200 165.200 ;
        RECT 12.700 165.100 13.000 165.800 ;
        RECT 14.600 165.600 15.000 165.800 ;
        RECT 16.600 165.400 17.200 165.800 ;
        RECT 18.200 165.400 18.600 166.200 ;
        RECT 19.000 166.100 19.300 166.800 ;
        RECT 20.600 166.100 21.000 166.600 ;
        RECT 19.000 165.800 21.000 166.100 ;
        RECT 21.400 165.800 21.700 167.300 ;
        RECT 23.000 167.400 24.900 167.700 ;
        RECT 16.600 165.100 16.900 165.400 ;
        RECT 19.000 165.100 19.300 165.800 ;
        RECT 21.400 165.400 22.000 165.800 ;
        RECT 23.000 165.700 23.400 167.400 ;
        RECT 26.500 167.100 26.900 167.200 ;
        RECT 29.400 167.100 29.700 168.200 ;
        RECT 31.800 167.500 32.200 169.900 ;
        RECT 32.600 167.700 33.000 169.900 ;
        RECT 34.700 169.200 35.300 169.900 ;
        RECT 34.700 168.900 35.400 169.200 ;
        RECT 37.000 168.900 37.400 169.900 ;
        RECT 39.200 169.200 39.600 169.900 ;
        RECT 39.200 168.900 40.200 169.200 ;
        RECT 35.000 168.500 35.400 168.900 ;
        RECT 37.100 168.600 37.400 168.900 ;
        RECT 37.100 168.300 38.500 168.600 ;
        RECT 38.100 168.200 38.500 168.300 ;
        RECT 39.000 168.200 39.400 168.600 ;
        RECT 39.800 168.500 40.200 168.900 ;
        RECT 34.100 167.700 34.500 167.800 ;
        RECT 32.600 167.400 34.500 167.700 ;
        RECT 31.000 167.100 31.800 167.200 ;
        RECT 26.300 166.800 31.800 167.100 ;
        RECT 25.400 166.400 25.800 166.500 ;
        RECT 23.900 166.100 25.800 166.400 ;
        RECT 23.900 166.000 24.300 166.100 ;
        RECT 24.700 165.700 25.100 165.800 ;
        RECT 23.000 165.400 25.100 165.700 ;
        RECT 21.400 165.100 21.700 165.400 ;
        RECT 10.700 164.800 11.200 165.100 ;
        RECT 11.500 164.800 12.200 165.100 ;
        RECT 10.700 161.100 11.100 164.800 ;
        RECT 11.500 164.200 11.800 164.800 ;
        RECT 11.400 163.800 11.800 164.200 ;
        RECT 12.600 161.100 13.000 165.100 ;
        RECT 13.400 164.800 15.400 165.100 ;
        RECT 13.400 161.100 13.800 164.800 ;
        RECT 15.000 161.100 15.400 164.800 ;
        RECT 15.800 164.800 16.900 165.100 ;
        RECT 15.800 161.100 16.200 164.800 ;
        RECT 18.500 164.700 19.400 165.100 ;
        RECT 20.600 164.800 21.700 165.100 ;
        RECT 18.500 161.100 18.900 164.700 ;
        RECT 20.600 161.100 21.000 164.800 ;
        RECT 23.000 161.100 23.400 165.400 ;
        RECT 26.300 165.200 26.600 166.800 ;
        RECT 29.900 166.700 30.300 166.800 ;
        RECT 29.400 166.200 29.800 166.300 ;
        RECT 30.700 166.200 31.100 166.300 ;
        RECT 28.600 165.900 31.100 166.200 ;
        RECT 28.600 165.800 29.000 165.900 ;
        RECT 32.600 165.700 33.000 167.400 ;
        RECT 36.100 167.100 36.500 167.200 ;
        RECT 39.000 167.100 39.300 168.200 ;
        RECT 41.400 167.500 41.800 169.900 ;
        RECT 43.000 168.900 43.400 169.900 ;
        RECT 42.200 167.800 42.600 168.600 ;
        RECT 43.100 167.200 43.400 168.900 ;
        RECT 40.600 167.100 41.400 167.200 ;
        RECT 35.900 166.800 41.400 167.100 ;
        RECT 43.000 166.800 43.400 167.200 ;
        RECT 46.200 168.500 46.600 169.500 ;
        RECT 46.200 167.400 46.500 168.500 ;
        RECT 48.300 168.000 48.700 169.500 ;
        RECT 48.300 167.700 49.100 168.000 ;
        RECT 48.700 167.500 49.100 167.700 ;
        RECT 46.200 167.100 48.300 167.400 ;
        RECT 35.000 166.400 35.400 166.500 ;
        RECT 33.500 166.100 35.400 166.400 ;
        RECT 33.500 166.000 33.900 166.100 ;
        RECT 34.300 165.700 34.700 165.800 ;
        RECT 29.400 165.500 32.200 165.600 ;
        RECT 29.300 165.400 32.200 165.500 ;
        RECT 25.400 164.900 26.600 165.200 ;
        RECT 27.300 165.300 32.200 165.400 ;
        RECT 27.300 165.100 29.700 165.300 ;
        RECT 25.400 164.400 25.700 164.900 ;
        RECT 25.000 164.000 25.700 164.400 ;
        RECT 26.500 164.500 26.900 164.600 ;
        RECT 27.300 164.500 27.600 165.100 ;
        RECT 26.500 164.200 27.600 164.500 ;
        RECT 27.900 164.500 30.600 164.800 ;
        RECT 27.900 164.400 28.300 164.500 ;
        RECT 30.200 164.400 30.600 164.500 ;
        RECT 27.100 163.700 27.500 163.800 ;
        RECT 28.500 163.700 28.900 163.800 ;
        RECT 25.400 163.100 25.800 163.500 ;
        RECT 27.100 163.400 28.900 163.700 ;
        RECT 27.500 163.100 27.800 163.400 ;
        RECT 30.200 163.100 30.600 163.500 ;
        RECT 25.100 161.100 25.700 163.100 ;
        RECT 27.400 161.100 27.800 163.100 ;
        RECT 29.600 162.800 30.600 163.100 ;
        RECT 29.600 161.100 30.000 162.800 ;
        RECT 31.800 161.100 32.200 165.300 ;
        RECT 32.600 165.400 34.700 165.700 ;
        RECT 32.600 161.100 33.000 165.400 ;
        RECT 35.900 165.200 36.200 166.800 ;
        RECT 39.500 166.700 39.900 166.800 ;
        RECT 39.000 166.200 39.400 166.300 ;
        RECT 40.300 166.200 40.700 166.300 ;
        RECT 43.100 166.200 43.400 166.800 ;
        RECT 47.800 166.900 48.300 167.100 ;
        RECT 48.800 167.200 49.100 167.500 ;
        RECT 51.000 167.700 51.400 169.900 ;
        RECT 53.100 169.200 53.700 169.900 ;
        RECT 53.100 168.900 53.800 169.200 ;
        RECT 55.400 168.900 55.800 169.900 ;
        RECT 57.600 169.200 58.000 169.900 ;
        RECT 57.600 168.900 58.600 169.200 ;
        RECT 53.400 168.500 53.800 168.900 ;
        RECT 55.500 168.600 55.800 168.900 ;
        RECT 55.500 168.300 56.900 168.600 ;
        RECT 56.500 168.200 56.900 168.300 ;
        RECT 57.400 168.200 57.800 168.600 ;
        RECT 58.200 168.500 58.600 168.900 ;
        RECT 52.500 167.700 52.900 167.800 ;
        RECT 51.000 167.400 52.900 167.700 ;
        RECT 38.200 165.900 40.700 166.200 ;
        RECT 38.200 165.800 38.600 165.900 ;
        RECT 43.000 165.800 43.400 166.200 ;
        RECT 39.000 165.500 41.800 165.600 ;
        RECT 38.900 165.400 41.800 165.500 ;
        RECT 35.000 164.900 36.200 165.200 ;
        RECT 36.900 165.300 41.800 165.400 ;
        RECT 36.900 165.100 39.300 165.300 ;
        RECT 35.000 164.400 35.300 164.900 ;
        RECT 34.600 164.000 35.300 164.400 ;
        RECT 36.100 164.500 36.500 164.600 ;
        RECT 36.900 164.500 37.200 165.100 ;
        RECT 36.100 164.200 37.200 164.500 ;
        RECT 37.500 164.500 40.200 164.800 ;
        RECT 37.500 164.400 37.900 164.500 ;
        RECT 39.800 164.400 40.200 164.500 ;
        RECT 36.700 163.700 37.100 163.800 ;
        RECT 38.100 163.700 38.500 163.800 ;
        RECT 35.000 163.100 35.400 163.500 ;
        RECT 36.700 163.400 38.500 163.700 ;
        RECT 37.100 163.100 37.400 163.400 ;
        RECT 39.800 163.100 40.200 163.500 ;
        RECT 34.700 161.100 35.300 163.100 ;
        RECT 37.000 161.100 37.400 163.100 ;
        RECT 39.200 162.800 40.200 163.100 ;
        RECT 39.200 161.100 39.600 162.800 ;
        RECT 41.400 161.100 41.800 165.300 ;
        RECT 43.100 165.100 43.400 165.800 ;
        RECT 43.800 165.400 44.200 166.200 ;
        RECT 44.600 166.100 45.000 166.200 ;
        RECT 46.200 166.100 46.600 166.600 ;
        RECT 44.600 165.800 46.600 166.100 ;
        RECT 47.000 165.800 47.400 166.600 ;
        RECT 47.800 166.500 48.500 166.900 ;
        RECT 48.800 166.800 49.800 167.200 ;
        RECT 47.800 165.500 48.100 166.500 ;
        RECT 48.800 166.200 49.100 166.800 ;
        RECT 48.600 165.800 49.100 166.200 ;
        RECT 46.200 165.200 48.100 165.500 ;
        RECT 43.000 164.700 43.900 165.100 ;
        RECT 43.500 161.100 43.900 164.700 ;
        RECT 46.200 163.500 46.500 165.200 ;
        RECT 48.800 164.900 49.100 165.800 ;
        RECT 49.400 165.400 49.800 166.200 ;
        RECT 51.000 165.700 51.400 167.400 ;
        RECT 54.500 167.100 54.900 167.200 ;
        RECT 57.400 167.100 57.700 168.200 ;
        RECT 59.800 167.500 60.200 169.900 ;
        RECT 61.400 168.900 61.800 169.900 ;
        RECT 61.400 167.200 61.700 168.900 ;
        RECT 62.200 167.800 62.600 168.600 ;
        RECT 63.000 167.700 63.400 169.900 ;
        RECT 65.100 169.200 65.700 169.900 ;
        RECT 65.100 168.900 65.800 169.200 ;
        RECT 67.400 168.900 67.800 169.900 ;
        RECT 69.600 169.200 70.000 169.900 ;
        RECT 69.600 168.900 70.600 169.200 ;
        RECT 65.400 168.500 65.800 168.900 ;
        RECT 67.500 168.600 67.800 168.900 ;
        RECT 67.500 168.300 68.900 168.600 ;
        RECT 68.500 168.200 68.900 168.300 ;
        RECT 69.400 168.200 69.800 168.600 ;
        RECT 70.200 168.500 70.600 168.900 ;
        RECT 64.500 167.700 64.900 167.800 ;
        RECT 63.000 167.400 64.900 167.700 ;
        RECT 59.000 167.100 59.800 167.200 ;
        RECT 54.300 166.800 59.800 167.100 ;
        RECT 61.400 166.800 61.800 167.200 ;
        RECT 53.400 166.400 53.800 166.500 ;
        RECT 51.900 166.100 53.800 166.400 ;
        RECT 54.300 166.100 54.600 166.800 ;
        RECT 57.900 166.700 58.300 166.800 ;
        RECT 57.400 166.200 57.800 166.300 ;
        RECT 58.700 166.200 59.100 166.300 ;
        RECT 55.000 166.100 55.400 166.200 ;
        RECT 51.900 166.000 52.300 166.100 ;
        RECT 54.200 165.800 55.400 166.100 ;
        RECT 56.600 165.900 59.100 166.200 ;
        RECT 56.600 165.800 57.000 165.900 ;
        RECT 52.700 165.700 53.100 165.800 ;
        RECT 51.000 165.400 53.100 165.700 ;
        RECT 48.300 164.600 49.100 164.900 ;
        RECT 46.200 161.500 46.600 163.500 ;
        RECT 48.300 161.100 48.700 164.600 ;
        RECT 51.000 161.100 51.400 165.400 ;
        RECT 54.300 165.200 54.600 165.800 ;
        RECT 57.400 165.500 60.200 165.600 ;
        RECT 57.300 165.400 60.200 165.500 ;
        RECT 60.600 165.400 61.000 166.200 ;
        RECT 61.400 166.100 61.700 166.800 ;
        RECT 62.200 166.100 62.600 166.200 ;
        RECT 61.400 165.800 62.600 166.100 ;
        RECT 53.400 164.900 54.600 165.200 ;
        RECT 55.300 165.300 60.200 165.400 ;
        RECT 55.300 165.100 57.700 165.300 ;
        RECT 53.400 164.400 53.700 164.900 ;
        RECT 53.000 164.000 53.700 164.400 ;
        RECT 54.500 164.500 54.900 164.600 ;
        RECT 55.300 164.500 55.600 165.100 ;
        RECT 54.500 164.200 55.600 164.500 ;
        RECT 55.900 164.500 58.600 164.800 ;
        RECT 55.900 164.400 56.300 164.500 ;
        RECT 58.200 164.400 58.600 164.500 ;
        RECT 55.100 163.700 55.500 163.800 ;
        RECT 56.500 163.700 56.900 163.800 ;
        RECT 53.400 163.100 53.800 163.500 ;
        RECT 55.100 163.400 56.900 163.700 ;
        RECT 55.500 163.100 55.800 163.400 ;
        RECT 58.200 163.100 58.600 163.500 ;
        RECT 53.100 161.100 53.700 163.100 ;
        RECT 55.400 161.100 55.800 163.100 ;
        RECT 57.600 162.800 58.600 163.100 ;
        RECT 57.600 161.100 58.000 162.800 ;
        RECT 59.800 161.100 60.200 165.300 ;
        RECT 61.400 165.100 61.700 165.800 ;
        RECT 63.000 165.700 63.400 167.400 ;
        RECT 69.400 167.200 69.700 168.200 ;
        RECT 71.800 167.500 72.200 169.900 ;
        RECT 72.600 167.700 73.000 169.900 ;
        RECT 74.700 169.200 75.300 169.900 ;
        RECT 74.700 168.900 75.400 169.200 ;
        RECT 77.000 168.900 77.400 169.900 ;
        RECT 79.200 169.200 79.600 169.900 ;
        RECT 79.200 168.900 80.200 169.200 ;
        RECT 75.000 168.500 75.400 168.900 ;
        RECT 77.100 168.600 77.400 168.900 ;
        RECT 77.100 168.300 78.500 168.600 ;
        RECT 78.100 168.200 78.500 168.300 ;
        RECT 79.000 168.200 79.400 168.600 ;
        RECT 79.800 168.500 80.200 168.900 ;
        RECT 74.100 167.700 74.500 167.800 ;
        RECT 72.600 167.400 74.500 167.700 ;
        RECT 66.500 167.100 66.900 167.200 ;
        RECT 69.400 167.100 69.800 167.200 ;
        RECT 71.000 167.100 71.800 167.200 ;
        RECT 66.300 166.800 71.800 167.100 ;
        RECT 65.400 166.400 65.800 166.500 ;
        RECT 63.900 166.100 65.800 166.400 ;
        RECT 63.900 166.000 64.300 166.100 ;
        RECT 64.700 165.700 65.100 165.800 ;
        RECT 63.000 165.400 65.100 165.700 ;
        RECT 60.900 164.700 61.800 165.100 ;
        RECT 60.900 161.100 61.300 164.700 ;
        RECT 63.000 161.100 63.400 165.400 ;
        RECT 66.300 165.200 66.600 166.800 ;
        RECT 69.900 166.700 70.300 166.800 ;
        RECT 70.700 166.200 71.100 166.300 ;
        RECT 67.000 166.100 67.400 166.200 ;
        RECT 68.600 166.100 71.100 166.200 ;
        RECT 67.000 165.900 71.100 166.100 ;
        RECT 67.000 165.800 69.000 165.900 ;
        RECT 72.600 165.700 73.000 167.400 ;
        RECT 76.100 167.100 76.500 167.200 ;
        RECT 79.000 167.100 79.300 168.200 ;
        RECT 81.400 167.500 81.800 169.900 ;
        RECT 83.800 167.600 84.200 169.900 ;
        RECT 85.400 168.900 85.800 169.900 ;
        RECT 84.600 167.800 85.000 168.600 ;
        RECT 83.100 167.300 84.200 167.600 ;
        RECT 80.600 167.100 81.400 167.200 ;
        RECT 75.900 166.800 81.400 167.100 ;
        RECT 75.000 166.400 75.400 166.500 ;
        RECT 73.500 166.100 75.400 166.400 ;
        RECT 73.500 166.000 73.900 166.100 ;
        RECT 74.300 165.700 74.700 165.800 ;
        RECT 69.400 165.500 72.200 165.600 ;
        RECT 69.300 165.400 72.200 165.500 ;
        RECT 65.400 164.900 66.600 165.200 ;
        RECT 67.300 165.300 72.200 165.400 ;
        RECT 67.300 165.100 69.700 165.300 ;
        RECT 65.400 164.400 65.700 164.900 ;
        RECT 65.000 164.000 65.700 164.400 ;
        RECT 66.500 164.500 66.900 164.600 ;
        RECT 67.300 164.500 67.600 165.100 ;
        RECT 66.500 164.200 67.600 164.500 ;
        RECT 67.900 164.500 70.600 164.800 ;
        RECT 67.900 164.400 68.300 164.500 ;
        RECT 70.200 164.400 70.600 164.500 ;
        RECT 67.100 163.700 67.500 163.800 ;
        RECT 68.500 163.700 68.900 163.800 ;
        RECT 65.400 163.100 65.800 163.500 ;
        RECT 67.100 163.400 68.900 163.700 ;
        RECT 67.500 163.100 67.800 163.400 ;
        RECT 70.200 163.100 70.600 163.500 ;
        RECT 65.100 161.100 65.700 163.100 ;
        RECT 67.400 161.100 67.800 163.100 ;
        RECT 69.600 162.800 70.600 163.100 ;
        RECT 69.600 161.100 70.000 162.800 ;
        RECT 71.800 161.100 72.200 165.300 ;
        RECT 72.600 165.400 74.700 165.700 ;
        RECT 72.600 161.100 73.000 165.400 ;
        RECT 75.900 165.200 76.200 166.800 ;
        RECT 79.500 166.700 79.900 166.800 ;
        RECT 79.000 166.200 79.400 166.300 ;
        RECT 80.300 166.200 80.700 166.300 ;
        RECT 78.200 165.900 80.700 166.200 ;
        RECT 78.200 165.800 78.600 165.900 ;
        RECT 83.100 165.800 83.400 167.300 ;
        RECT 85.500 167.200 85.800 168.900 ;
        RECT 88.600 167.600 89.000 169.900 ;
        RECT 85.400 166.800 85.800 167.200 ;
        RECT 83.800 166.100 84.200 166.600 ;
        RECT 85.500 166.100 85.800 166.800 ;
        RECT 87.900 167.300 89.000 167.600 ;
        RECT 83.800 165.800 85.800 166.100 ;
        RECT 79.000 165.500 81.800 165.600 ;
        RECT 78.900 165.400 81.800 165.500 ;
        RECT 82.800 165.400 83.400 165.800 ;
        RECT 75.000 164.900 76.200 165.200 ;
        RECT 76.900 165.300 81.800 165.400 ;
        RECT 76.900 165.100 79.300 165.300 ;
        RECT 75.000 164.400 75.300 164.900 ;
        RECT 74.600 164.000 75.300 164.400 ;
        RECT 76.100 164.500 76.500 164.600 ;
        RECT 76.900 164.500 77.200 165.100 ;
        RECT 76.100 164.200 77.200 164.500 ;
        RECT 77.500 164.500 80.200 164.800 ;
        RECT 77.500 164.400 77.900 164.500 ;
        RECT 79.800 164.400 80.200 164.500 ;
        RECT 76.700 163.700 77.100 163.800 ;
        RECT 78.100 163.700 78.500 163.800 ;
        RECT 75.000 163.100 75.400 163.500 ;
        RECT 76.700 163.400 78.500 163.700 ;
        RECT 77.100 163.100 77.400 163.400 ;
        RECT 79.800 163.100 80.200 163.500 ;
        RECT 74.700 161.100 75.300 163.100 ;
        RECT 77.000 161.100 77.400 163.100 ;
        RECT 79.200 162.800 80.200 163.100 ;
        RECT 79.200 161.100 79.600 162.800 ;
        RECT 81.400 161.100 81.800 165.300 ;
        RECT 83.100 165.100 83.400 165.400 ;
        RECT 85.500 165.100 85.800 165.800 ;
        RECT 86.200 165.400 86.600 166.200 ;
        RECT 87.900 165.800 88.200 167.300 ;
        RECT 88.600 166.100 89.000 166.600 ;
        RECT 89.400 166.100 89.800 169.900 ;
        RECT 90.200 167.800 90.600 168.600 ;
        RECT 88.600 165.800 89.800 166.100 ;
        RECT 87.600 165.400 88.200 165.800 ;
        RECT 87.900 165.100 88.200 165.400 ;
        RECT 83.100 164.800 84.200 165.100 ;
        RECT 83.800 161.100 84.200 164.800 ;
        RECT 85.400 164.700 86.300 165.100 ;
        RECT 87.900 164.800 89.000 165.100 ;
        RECT 85.900 161.100 86.300 164.700 ;
        RECT 88.600 161.100 89.000 164.800 ;
        RECT 89.400 161.100 89.800 165.800 ;
        RECT 91.000 167.700 91.400 169.900 ;
        RECT 93.100 169.200 93.700 169.900 ;
        RECT 93.100 168.900 93.800 169.200 ;
        RECT 95.400 168.900 95.800 169.900 ;
        RECT 97.600 169.200 98.000 169.900 ;
        RECT 97.600 168.900 98.600 169.200 ;
        RECT 93.400 168.500 93.800 168.900 ;
        RECT 95.500 168.600 95.800 168.900 ;
        RECT 95.500 168.300 96.900 168.600 ;
        RECT 96.500 168.200 96.900 168.300 ;
        RECT 97.400 168.200 97.800 168.600 ;
        RECT 98.200 168.500 98.600 168.900 ;
        RECT 92.500 167.700 92.900 167.800 ;
        RECT 91.000 167.400 92.900 167.700 ;
        RECT 91.000 165.700 91.400 167.400 ;
        RECT 94.500 167.100 94.900 167.200 ;
        RECT 97.400 167.100 97.700 168.200 ;
        RECT 99.800 167.500 100.200 169.900 ;
        RECT 103.000 168.900 103.400 169.900 ;
        RECT 102.200 167.800 102.600 168.600 ;
        RECT 103.100 167.200 103.400 168.900 ;
        RECT 104.600 167.600 105.000 169.900 ;
        RECT 107.000 167.700 107.400 169.900 ;
        RECT 109.100 169.200 109.700 169.900 ;
        RECT 109.100 168.900 109.800 169.200 ;
        RECT 111.400 168.900 111.800 169.900 ;
        RECT 113.600 169.200 114.000 169.900 ;
        RECT 113.600 168.900 114.600 169.200 ;
        RECT 109.400 168.500 109.800 168.900 ;
        RECT 111.500 168.600 111.800 168.900 ;
        RECT 111.500 168.300 112.900 168.600 ;
        RECT 112.500 168.200 112.900 168.300 ;
        RECT 113.400 168.200 113.800 168.600 ;
        RECT 114.200 168.500 114.600 168.900 ;
        RECT 108.500 167.700 108.900 167.800 ;
        RECT 104.600 167.300 105.700 167.600 ;
        RECT 99.000 167.100 99.800 167.200 ;
        RECT 94.300 166.800 99.800 167.100 ;
        RECT 103.000 166.800 103.400 167.200 ;
        RECT 93.400 166.400 93.800 166.500 ;
        RECT 91.900 166.100 93.800 166.400 ;
        RECT 94.300 166.200 94.600 166.800 ;
        RECT 97.900 166.700 98.300 166.800 ;
        RECT 97.400 166.200 97.800 166.300 ;
        RECT 98.700 166.200 99.100 166.300 ;
        RECT 91.900 166.000 92.300 166.100 ;
        RECT 94.200 165.800 94.600 166.200 ;
        RECT 96.600 165.900 99.100 166.200 ;
        RECT 101.400 166.100 101.800 166.200 ;
        RECT 103.100 166.100 103.400 166.800 ;
        RECT 96.600 165.800 97.000 165.900 ;
        RECT 101.400 165.800 103.400 166.100 ;
        RECT 92.700 165.700 93.100 165.800 ;
        RECT 91.000 165.400 93.100 165.700 ;
        RECT 91.000 161.100 91.400 165.400 ;
        RECT 94.300 165.200 94.600 165.800 ;
        RECT 97.400 165.500 100.200 165.600 ;
        RECT 97.300 165.400 100.200 165.500 ;
        RECT 93.400 164.900 94.600 165.200 ;
        RECT 95.300 165.300 100.200 165.400 ;
        RECT 95.300 165.100 97.700 165.300 ;
        RECT 93.400 164.400 93.700 164.900 ;
        RECT 93.000 164.000 93.700 164.400 ;
        RECT 94.500 164.500 94.900 164.600 ;
        RECT 95.300 164.500 95.600 165.100 ;
        RECT 94.500 164.200 95.600 164.500 ;
        RECT 95.900 164.500 98.600 164.800 ;
        RECT 95.900 164.400 96.300 164.500 ;
        RECT 98.200 164.400 98.600 164.500 ;
        RECT 95.100 163.700 95.500 163.800 ;
        RECT 96.500 163.700 96.900 163.800 ;
        RECT 93.400 163.100 93.800 163.500 ;
        RECT 95.100 163.400 96.900 163.700 ;
        RECT 95.500 163.100 95.800 163.400 ;
        RECT 98.200 163.100 98.600 163.500 ;
        RECT 93.100 161.100 93.700 163.100 ;
        RECT 95.400 161.100 95.800 163.100 ;
        RECT 97.600 162.800 98.600 163.100 ;
        RECT 97.600 161.100 98.000 162.800 ;
        RECT 99.800 161.100 100.200 165.300 ;
        RECT 103.100 165.100 103.400 165.800 ;
        RECT 103.800 165.400 104.200 166.200 ;
        RECT 105.400 165.800 105.700 167.300 ;
        RECT 107.000 167.400 108.900 167.700 ;
        RECT 105.400 165.400 106.000 165.800 ;
        RECT 107.000 165.700 107.400 167.400 ;
        RECT 110.500 167.100 110.900 167.200 ;
        RECT 113.400 167.100 113.700 168.200 ;
        RECT 115.800 167.500 116.200 169.900 ;
        RECT 118.200 167.600 118.600 169.900 ;
        RECT 117.500 167.300 118.600 167.600 ;
        RECT 119.000 167.600 119.400 169.900 ;
        RECT 121.400 167.700 121.800 169.900 ;
        RECT 123.500 169.200 124.100 169.900 ;
        RECT 123.500 168.900 124.200 169.200 ;
        RECT 125.800 168.900 126.200 169.900 ;
        RECT 128.000 169.200 128.400 169.900 ;
        RECT 128.000 168.900 129.000 169.200 ;
        RECT 123.800 168.500 124.200 168.900 ;
        RECT 125.900 168.600 126.200 168.900 ;
        RECT 125.900 168.300 127.300 168.600 ;
        RECT 126.900 168.200 127.300 168.300 ;
        RECT 127.800 168.200 128.200 168.600 ;
        RECT 128.600 168.500 129.000 168.900 ;
        RECT 122.900 167.700 123.300 167.800 ;
        RECT 119.000 167.300 120.100 167.600 ;
        RECT 115.000 167.100 115.800 167.200 ;
        RECT 110.300 166.800 115.800 167.100 ;
        RECT 109.400 166.400 109.800 166.500 ;
        RECT 107.900 166.100 109.800 166.400 ;
        RECT 107.900 166.000 108.300 166.100 ;
        RECT 108.700 165.700 109.100 165.800 ;
        RECT 107.000 165.400 109.100 165.700 ;
        RECT 105.400 165.100 105.700 165.400 ;
        RECT 103.000 164.700 103.900 165.100 ;
        RECT 103.500 161.100 103.900 164.700 ;
        RECT 104.600 164.800 105.700 165.100 ;
        RECT 104.600 161.100 105.000 164.800 ;
        RECT 107.000 161.100 107.400 165.400 ;
        RECT 110.300 165.200 110.600 166.800 ;
        RECT 113.900 166.700 114.300 166.800 ;
        RECT 114.700 166.200 115.100 166.300 ;
        RECT 112.600 165.900 115.100 166.200 ;
        RECT 112.600 165.800 113.000 165.900 ;
        RECT 117.500 165.800 117.800 167.300 ;
        RECT 118.200 165.800 118.600 166.600 ;
        RECT 119.000 165.800 119.400 166.600 ;
        RECT 119.800 165.800 120.100 167.300 ;
        RECT 121.400 167.400 123.300 167.700 ;
        RECT 113.400 165.500 116.200 165.600 ;
        RECT 113.300 165.400 116.200 165.500 ;
        RECT 117.200 165.400 117.800 165.800 ;
        RECT 109.400 164.900 110.600 165.200 ;
        RECT 111.300 165.300 116.200 165.400 ;
        RECT 111.300 165.100 113.700 165.300 ;
        RECT 109.400 164.400 109.700 164.900 ;
        RECT 109.000 164.000 109.700 164.400 ;
        RECT 110.500 164.500 110.900 164.600 ;
        RECT 111.300 164.500 111.600 165.100 ;
        RECT 110.500 164.200 111.600 164.500 ;
        RECT 111.900 164.500 114.600 164.800 ;
        RECT 111.900 164.400 112.300 164.500 ;
        RECT 114.200 164.400 114.600 164.500 ;
        RECT 111.100 163.700 111.500 163.800 ;
        RECT 112.500 163.700 112.900 163.800 ;
        RECT 109.400 163.100 109.800 163.500 ;
        RECT 111.100 163.400 112.900 163.700 ;
        RECT 111.500 163.100 111.800 163.400 ;
        RECT 114.200 163.100 114.600 163.500 ;
        RECT 109.100 161.100 109.700 163.100 ;
        RECT 111.400 161.100 111.800 163.100 ;
        RECT 113.600 162.800 114.600 163.100 ;
        RECT 113.600 161.100 114.000 162.800 ;
        RECT 115.800 161.100 116.200 165.300 ;
        RECT 117.500 165.100 117.800 165.400 ;
        RECT 119.800 165.400 120.400 165.800 ;
        RECT 121.400 165.700 121.800 167.400 ;
        RECT 124.900 167.100 125.300 167.200 ;
        RECT 127.800 167.100 128.100 168.200 ;
        RECT 130.200 167.500 130.600 169.900 ;
        RECT 132.600 167.600 133.000 169.900 ;
        RECT 131.900 167.300 133.000 167.600 ;
        RECT 133.400 167.600 133.800 169.900 ;
        RECT 133.400 167.300 134.500 167.600 ;
        RECT 135.800 167.500 136.200 169.900 ;
        RECT 138.000 169.200 138.400 169.900 ;
        RECT 137.400 168.900 138.400 169.200 ;
        RECT 140.200 168.900 140.600 169.900 ;
        RECT 142.300 169.200 142.900 169.900 ;
        RECT 142.200 168.900 142.900 169.200 ;
        RECT 137.400 168.500 137.800 168.900 ;
        RECT 140.200 168.600 140.500 168.900 ;
        RECT 138.200 168.200 138.600 168.600 ;
        RECT 139.100 168.300 140.500 168.600 ;
        RECT 142.200 168.500 142.600 168.900 ;
        RECT 139.100 168.200 139.500 168.300 ;
        RECT 129.400 167.100 130.200 167.200 ;
        RECT 124.700 166.800 130.200 167.100 ;
        RECT 123.800 166.400 124.200 166.500 ;
        RECT 122.300 166.100 124.200 166.400 ;
        RECT 124.700 166.200 125.000 166.800 ;
        RECT 128.300 166.700 128.700 166.800 ;
        RECT 129.100 166.200 129.500 166.300 ;
        RECT 122.300 166.000 122.700 166.100 ;
        RECT 124.600 165.800 125.000 166.200 ;
        RECT 127.000 165.900 129.500 166.200 ;
        RECT 127.000 165.800 127.400 165.900 ;
        RECT 131.900 165.800 132.200 167.300 ;
        RECT 123.100 165.700 123.500 165.800 ;
        RECT 121.400 165.400 123.500 165.700 ;
        RECT 119.800 165.100 120.100 165.400 ;
        RECT 117.500 164.800 118.600 165.100 ;
        RECT 118.200 161.100 118.600 164.800 ;
        RECT 119.000 164.800 120.100 165.100 ;
        RECT 119.000 161.100 119.400 164.800 ;
        RECT 121.400 161.100 121.800 165.400 ;
        RECT 124.700 165.200 125.000 165.800 ;
        RECT 127.800 165.500 130.600 165.600 ;
        RECT 127.700 165.400 130.600 165.500 ;
        RECT 131.600 165.400 132.200 165.800 ;
        RECT 123.800 164.900 125.000 165.200 ;
        RECT 125.700 165.300 130.600 165.400 ;
        RECT 125.700 165.100 128.100 165.300 ;
        RECT 123.800 164.400 124.100 164.900 ;
        RECT 123.400 164.000 124.100 164.400 ;
        RECT 124.900 164.500 125.300 164.600 ;
        RECT 125.700 164.500 126.000 165.100 ;
        RECT 124.900 164.200 126.000 164.500 ;
        RECT 126.300 164.500 129.000 164.800 ;
        RECT 126.300 164.400 126.700 164.500 ;
        RECT 128.600 164.400 129.000 164.500 ;
        RECT 125.500 163.700 125.900 163.800 ;
        RECT 126.900 163.700 127.300 163.800 ;
        RECT 123.800 163.100 124.200 163.500 ;
        RECT 125.500 163.400 127.300 163.700 ;
        RECT 125.900 163.100 126.200 163.400 ;
        RECT 128.600 163.100 129.000 163.500 ;
        RECT 123.500 161.100 124.100 163.100 ;
        RECT 125.800 161.100 126.200 163.100 ;
        RECT 128.000 162.800 129.000 163.100 ;
        RECT 128.000 161.100 128.400 162.800 ;
        RECT 130.200 161.100 130.600 165.300 ;
        RECT 131.900 165.100 132.200 165.400 ;
        RECT 134.200 165.800 134.500 167.300 ;
        RECT 138.300 167.200 138.600 168.200 ;
        RECT 143.100 167.700 143.500 167.800 ;
        RECT 144.600 167.700 145.000 169.900 ;
        RECT 146.200 168.900 146.600 169.900 ;
        RECT 145.400 167.800 145.800 168.600 ;
        RECT 143.100 167.400 145.000 167.700 ;
        RECT 136.200 167.100 137.000 167.200 ;
        RECT 138.200 167.100 138.600 167.200 ;
        RECT 141.100 167.100 141.500 167.200 ;
        RECT 136.200 166.800 141.700 167.100 ;
        RECT 137.700 166.700 138.100 166.800 ;
        RECT 136.900 166.200 137.300 166.300 ;
        RECT 136.900 165.900 139.400 166.200 ;
        RECT 139.000 165.800 139.400 165.900 ;
        RECT 134.200 165.400 134.800 165.800 ;
        RECT 135.800 165.500 138.600 165.600 ;
        RECT 135.800 165.400 138.700 165.500 ;
        RECT 134.200 165.100 134.500 165.400 ;
        RECT 131.900 164.800 133.000 165.100 ;
        RECT 132.600 161.100 133.000 164.800 ;
        RECT 133.400 164.800 134.500 165.100 ;
        RECT 135.800 165.300 140.700 165.400 ;
        RECT 133.400 161.100 133.800 164.800 ;
        RECT 135.800 161.100 136.200 165.300 ;
        RECT 138.300 165.100 140.700 165.300 ;
        RECT 137.400 164.500 140.100 164.800 ;
        RECT 137.400 164.400 137.800 164.500 ;
        RECT 139.700 164.400 140.100 164.500 ;
        RECT 140.400 164.500 140.700 165.100 ;
        RECT 141.400 165.200 141.700 166.800 ;
        RECT 142.200 166.400 142.600 166.500 ;
        RECT 142.200 166.100 144.100 166.400 ;
        RECT 143.700 166.000 144.100 166.100 ;
        RECT 142.900 165.700 143.300 165.800 ;
        RECT 144.600 165.700 145.000 167.400 ;
        RECT 146.300 167.200 146.600 168.900 ;
        RECT 146.200 167.100 146.600 167.200 ;
        RECT 149.400 168.500 149.800 169.500 ;
        RECT 149.400 167.400 149.700 168.500 ;
        RECT 151.500 168.200 151.900 169.500 ;
        RECT 151.000 168.000 151.900 168.200 ;
        RECT 151.000 167.800 152.300 168.000 ;
        RECT 151.500 167.700 152.300 167.800 ;
        RECT 151.900 167.500 152.300 167.700 ;
        RECT 149.400 167.100 151.500 167.400 ;
        RECT 145.400 166.800 146.600 167.100 ;
        RECT 145.400 166.200 145.700 166.800 ;
        RECT 145.400 165.800 145.800 166.200 ;
        RECT 142.900 165.400 145.000 165.700 ;
        RECT 141.400 164.900 142.600 165.200 ;
        RECT 141.100 164.500 141.500 164.600 ;
        RECT 140.400 164.200 141.500 164.500 ;
        RECT 142.300 164.400 142.600 164.900 ;
        RECT 142.300 164.000 143.000 164.400 ;
        RECT 139.100 163.700 139.500 163.800 ;
        RECT 140.500 163.700 140.900 163.800 ;
        RECT 137.400 163.100 137.800 163.500 ;
        RECT 139.100 163.400 140.900 163.700 ;
        RECT 140.200 163.100 140.500 163.400 ;
        RECT 142.200 163.100 142.600 163.500 ;
        RECT 137.400 162.800 138.400 163.100 ;
        RECT 138.000 161.100 138.400 162.800 ;
        RECT 140.200 161.100 140.600 163.100 ;
        RECT 142.300 161.100 142.900 163.100 ;
        RECT 144.600 161.100 145.000 165.400 ;
        RECT 146.300 165.100 146.600 166.800 ;
        RECT 151.000 166.900 151.500 167.100 ;
        RECT 152.000 167.200 152.300 167.500 ;
        RECT 154.200 167.700 154.600 169.900 ;
        RECT 156.300 169.200 156.900 169.900 ;
        RECT 156.300 168.900 157.000 169.200 ;
        RECT 158.600 168.900 159.000 169.900 ;
        RECT 160.800 169.200 161.200 169.900 ;
        RECT 160.800 168.900 161.800 169.200 ;
        RECT 156.600 168.500 157.000 168.900 ;
        RECT 158.700 168.600 159.000 168.900 ;
        RECT 158.700 168.300 160.100 168.600 ;
        RECT 159.700 168.200 160.100 168.300 ;
        RECT 160.600 168.200 161.000 168.600 ;
        RECT 161.400 168.500 161.800 168.900 ;
        RECT 155.700 167.700 156.100 167.800 ;
        RECT 154.200 167.400 156.100 167.700 ;
        RECT 147.000 165.400 147.400 166.200 ;
        RECT 149.400 165.800 149.800 166.600 ;
        RECT 150.200 165.800 150.600 166.600 ;
        RECT 151.000 166.500 151.700 166.900 ;
        RECT 152.000 166.800 153.000 167.200 ;
        RECT 151.000 165.500 151.300 166.500 ;
        RECT 149.400 165.200 151.300 165.500 ;
        RECT 146.200 164.700 147.100 165.100 ;
        RECT 146.700 161.100 147.100 164.700 ;
        RECT 149.400 163.500 149.700 165.200 ;
        RECT 152.000 164.900 152.300 166.800 ;
        RECT 151.500 164.600 152.300 164.900 ;
        RECT 154.200 165.700 154.600 167.400 ;
        RECT 160.600 167.200 160.900 168.200 ;
        RECT 163.000 167.500 163.400 169.900 ;
        RECT 163.800 167.500 164.200 169.900 ;
        RECT 166.000 169.200 166.400 169.900 ;
        RECT 165.400 168.900 166.400 169.200 ;
        RECT 168.200 168.900 168.600 169.900 ;
        RECT 170.300 169.200 170.900 169.900 ;
        RECT 170.200 168.900 170.900 169.200 ;
        RECT 165.400 168.500 165.800 168.900 ;
        RECT 168.200 168.600 168.500 168.900 ;
        RECT 166.200 168.200 166.600 168.600 ;
        RECT 167.100 168.300 168.500 168.600 ;
        RECT 170.200 168.500 170.600 168.900 ;
        RECT 167.100 168.200 167.500 168.300 ;
        RECT 157.700 167.100 158.100 167.200 ;
        RECT 160.600 167.100 161.000 167.200 ;
        RECT 162.200 167.100 163.000 167.200 ;
        RECT 157.500 166.800 163.000 167.100 ;
        RECT 164.200 167.100 165.000 167.200 ;
        RECT 166.300 167.100 166.600 168.200 ;
        RECT 171.100 167.700 171.500 167.800 ;
        RECT 172.600 167.700 173.000 169.900 ;
        RECT 171.100 167.400 173.000 167.700 ;
        RECT 169.100 167.100 169.500 167.200 ;
        RECT 164.200 166.800 169.700 167.100 ;
        RECT 156.600 166.400 157.000 166.500 ;
        RECT 155.100 166.100 157.000 166.400 ;
        RECT 155.100 166.000 155.500 166.100 ;
        RECT 155.900 165.700 156.300 165.800 ;
        RECT 154.200 165.400 156.300 165.700 ;
        RECT 149.400 161.500 149.800 163.500 ;
        RECT 151.500 161.100 151.900 164.600 ;
        RECT 154.200 161.100 154.600 165.400 ;
        RECT 157.500 165.200 157.800 166.800 ;
        RECT 161.100 166.700 161.500 166.800 ;
        RECT 165.700 166.700 166.100 166.800 ;
        RECT 161.900 166.200 162.300 166.300 ;
        RECT 159.800 165.900 162.300 166.200 ;
        RECT 164.900 166.200 165.300 166.300 ;
        RECT 169.400 166.200 169.700 166.800 ;
        RECT 170.200 166.400 170.600 166.500 ;
        RECT 164.900 165.900 167.400 166.200 ;
        RECT 159.800 165.800 160.200 165.900 ;
        RECT 167.000 165.800 167.400 165.900 ;
        RECT 169.400 165.800 169.800 166.200 ;
        RECT 170.200 166.100 172.100 166.400 ;
        RECT 171.700 166.000 172.100 166.100 ;
        RECT 160.600 165.500 163.400 165.600 ;
        RECT 160.500 165.400 163.400 165.500 ;
        RECT 156.600 164.900 157.800 165.200 ;
        RECT 158.500 165.300 163.400 165.400 ;
        RECT 158.500 165.100 160.900 165.300 ;
        RECT 156.600 164.400 156.900 164.900 ;
        RECT 156.200 164.000 156.900 164.400 ;
        RECT 157.700 164.500 158.100 164.600 ;
        RECT 158.500 164.500 158.800 165.100 ;
        RECT 157.700 164.200 158.800 164.500 ;
        RECT 159.100 164.500 161.800 164.800 ;
        RECT 159.100 164.400 159.500 164.500 ;
        RECT 161.400 164.400 161.800 164.500 ;
        RECT 158.300 163.700 158.700 163.800 ;
        RECT 159.700 163.700 160.100 163.800 ;
        RECT 156.600 163.100 157.000 163.500 ;
        RECT 158.300 163.400 160.100 163.700 ;
        RECT 158.700 163.100 159.000 163.400 ;
        RECT 161.400 163.100 161.800 163.500 ;
        RECT 156.300 161.100 156.900 163.100 ;
        RECT 158.600 161.100 159.000 163.100 ;
        RECT 160.800 162.800 161.800 163.100 ;
        RECT 160.800 161.100 161.200 162.800 ;
        RECT 163.000 161.100 163.400 165.300 ;
        RECT 163.800 165.500 166.600 165.600 ;
        RECT 163.800 165.400 166.700 165.500 ;
        RECT 163.800 165.300 168.700 165.400 ;
        RECT 163.800 161.100 164.200 165.300 ;
        RECT 166.300 165.100 168.700 165.300 ;
        RECT 165.400 164.500 168.100 164.800 ;
        RECT 165.400 164.400 165.800 164.500 ;
        RECT 167.700 164.400 168.100 164.500 ;
        RECT 168.400 164.500 168.700 165.100 ;
        RECT 169.400 165.200 169.700 165.800 ;
        RECT 170.900 165.700 171.300 165.800 ;
        RECT 172.600 165.700 173.000 167.400 ;
        RECT 173.400 167.600 173.800 169.900 ;
        RECT 175.800 167.700 176.200 169.900 ;
        RECT 177.900 169.200 178.500 169.900 ;
        RECT 177.900 168.900 178.600 169.200 ;
        RECT 180.200 168.900 180.600 169.900 ;
        RECT 182.400 169.200 182.800 169.900 ;
        RECT 182.400 168.900 183.400 169.200 ;
        RECT 178.200 168.500 178.600 168.900 ;
        RECT 180.300 168.600 180.600 168.900 ;
        RECT 180.300 168.300 181.700 168.600 ;
        RECT 181.300 168.200 181.700 168.300 ;
        RECT 182.200 168.200 182.600 168.600 ;
        RECT 183.000 168.500 183.400 168.900 ;
        RECT 177.300 167.700 177.700 167.800 ;
        RECT 173.400 167.300 174.500 167.600 ;
        RECT 170.900 165.400 173.000 165.700 ;
        RECT 169.400 164.900 170.600 165.200 ;
        RECT 169.100 164.500 169.500 164.600 ;
        RECT 168.400 164.200 169.500 164.500 ;
        RECT 170.300 164.400 170.600 164.900 ;
        RECT 170.300 164.000 171.000 164.400 ;
        RECT 167.100 163.700 167.500 163.800 ;
        RECT 168.500 163.700 168.900 163.800 ;
        RECT 165.400 163.100 165.800 163.500 ;
        RECT 167.100 163.400 168.900 163.700 ;
        RECT 168.200 163.100 168.500 163.400 ;
        RECT 170.200 163.100 170.600 163.500 ;
        RECT 165.400 162.800 166.400 163.100 ;
        RECT 166.000 161.100 166.400 162.800 ;
        RECT 168.200 161.100 168.600 163.100 ;
        RECT 170.300 161.100 170.900 163.100 ;
        RECT 172.600 161.100 173.000 165.400 ;
        RECT 174.200 165.800 174.500 167.300 ;
        RECT 175.800 167.400 177.700 167.700 ;
        RECT 174.200 165.400 174.800 165.800 ;
        RECT 175.800 165.700 176.200 167.400 ;
        RECT 179.300 167.100 179.700 167.200 ;
        RECT 182.200 167.100 182.500 168.200 ;
        RECT 184.600 167.500 185.000 169.900 ;
        RECT 187.000 167.600 187.400 169.900 ;
        RECT 186.300 167.300 187.400 167.600 ;
        RECT 187.800 167.600 188.200 169.900 ;
        RECT 190.200 167.600 190.600 169.900 ;
        RECT 192.600 167.800 193.000 168.600 ;
        RECT 187.800 167.300 188.900 167.600 ;
        RECT 190.200 167.300 191.300 167.600 ;
        RECT 183.800 167.100 184.600 167.200 ;
        RECT 179.100 166.800 184.600 167.100 ;
        RECT 178.200 166.400 178.600 166.500 ;
        RECT 176.700 166.100 178.600 166.400 ;
        RECT 179.100 166.100 179.400 166.800 ;
        RECT 182.700 166.700 183.100 166.800 ;
        RECT 183.500 166.200 183.900 166.300 ;
        RECT 179.800 166.100 180.200 166.200 ;
        RECT 176.700 166.000 177.100 166.100 ;
        RECT 179.000 165.800 180.200 166.100 ;
        RECT 181.400 165.900 183.900 166.200 ;
        RECT 181.400 165.800 181.800 165.900 ;
        RECT 186.300 165.800 186.600 167.300 ;
        RECT 177.500 165.700 177.900 165.800 ;
        RECT 175.800 165.400 177.900 165.700 ;
        RECT 174.200 165.100 174.500 165.400 ;
        RECT 173.400 164.800 174.500 165.100 ;
        RECT 173.400 161.100 173.800 164.800 ;
        RECT 175.800 161.100 176.200 165.400 ;
        RECT 179.100 165.200 179.400 165.800 ;
        RECT 182.200 165.500 185.000 165.600 ;
        RECT 182.100 165.400 185.000 165.500 ;
        RECT 186.000 165.400 186.600 165.800 ;
        RECT 178.200 164.900 179.400 165.200 ;
        RECT 180.100 165.300 185.000 165.400 ;
        RECT 180.100 165.100 182.500 165.300 ;
        RECT 178.200 164.400 178.500 164.900 ;
        RECT 177.800 164.000 178.500 164.400 ;
        RECT 179.300 164.500 179.700 164.600 ;
        RECT 180.100 164.500 180.400 165.100 ;
        RECT 179.300 164.200 180.400 164.500 ;
        RECT 180.700 164.500 183.400 164.800 ;
        RECT 180.700 164.400 181.100 164.500 ;
        RECT 183.000 164.400 183.400 164.500 ;
        RECT 179.900 163.700 180.300 163.800 ;
        RECT 181.300 163.700 181.700 163.800 ;
        RECT 178.200 163.100 178.600 163.500 ;
        RECT 179.900 163.400 181.700 163.700 ;
        RECT 180.300 163.100 180.600 163.400 ;
        RECT 183.000 163.100 183.400 163.500 ;
        RECT 177.900 161.100 178.500 163.100 ;
        RECT 180.200 161.100 180.600 163.100 ;
        RECT 182.400 162.800 183.400 163.100 ;
        RECT 182.400 161.100 182.800 162.800 ;
        RECT 184.600 161.100 185.000 165.300 ;
        RECT 186.300 165.100 186.600 165.400 ;
        RECT 188.600 165.800 188.900 167.300 ;
        RECT 191.000 165.800 191.300 167.300 ;
        RECT 188.600 165.400 189.200 165.800 ;
        RECT 191.000 165.400 191.600 165.800 ;
        RECT 188.600 165.100 188.900 165.400 ;
        RECT 191.000 165.100 191.300 165.400 ;
        RECT 186.300 164.800 187.400 165.100 ;
        RECT 187.000 161.100 187.400 164.800 ;
        RECT 187.800 164.800 188.900 165.100 ;
        RECT 190.200 164.800 191.300 165.100 ;
        RECT 187.800 161.100 188.200 164.800 ;
        RECT 190.200 161.100 190.600 164.800 ;
        RECT 193.400 162.100 193.800 169.900 ;
        RECT 194.200 162.100 194.600 162.200 ;
        RECT 193.400 161.800 194.600 162.100 ;
        RECT 193.400 161.100 193.800 161.800 ;
        RECT 0.600 155.600 1.000 159.900 ;
        RECT 2.700 157.900 3.300 159.900 ;
        RECT 5.000 157.900 5.400 159.900 ;
        RECT 7.200 158.200 7.600 159.900 ;
        RECT 7.200 157.900 8.200 158.200 ;
        RECT 3.000 157.500 3.400 157.900 ;
        RECT 5.100 157.600 5.400 157.900 ;
        RECT 4.700 157.300 6.500 157.600 ;
        RECT 7.800 157.500 8.200 157.900 ;
        RECT 4.700 157.200 5.100 157.300 ;
        RECT 6.100 157.200 6.500 157.300 ;
        RECT 2.600 156.600 3.300 157.000 ;
        RECT 3.000 156.100 3.300 156.600 ;
        RECT 4.100 156.500 5.200 156.800 ;
        RECT 4.100 156.400 4.500 156.500 ;
        RECT 3.000 155.800 4.200 156.100 ;
        RECT 0.600 155.300 2.700 155.600 ;
        RECT 0.600 153.600 1.000 155.300 ;
        RECT 2.300 155.200 2.700 155.300 ;
        RECT 1.500 154.900 1.900 155.000 ;
        RECT 1.500 154.600 3.400 154.900 ;
        RECT 3.000 154.500 3.400 154.600 ;
        RECT 3.900 154.200 4.200 155.800 ;
        RECT 4.900 155.900 5.200 156.500 ;
        RECT 5.500 156.500 5.900 156.600 ;
        RECT 7.800 156.500 8.200 156.600 ;
        RECT 5.500 156.200 8.200 156.500 ;
        RECT 4.900 155.700 7.300 155.900 ;
        RECT 9.400 155.700 9.800 159.900 ;
        RECT 12.100 159.200 12.500 159.900 ;
        RECT 12.100 158.800 13.000 159.200 ;
        RECT 12.100 156.400 12.500 158.800 ;
        RECT 14.200 157.500 14.600 159.500 ;
        RECT 4.900 155.600 9.800 155.700 ;
        RECT 11.700 156.100 12.500 156.400 ;
        RECT 6.900 155.500 9.800 155.600 ;
        RECT 7.000 155.400 9.800 155.500 ;
        RECT 6.200 155.100 6.600 155.200 ;
        RECT 10.200 155.100 10.600 155.200 ;
        RECT 11.000 155.100 11.400 155.600 ;
        RECT 6.200 154.800 8.700 155.100 ;
        RECT 10.200 154.800 11.400 155.100 ;
        RECT 8.300 154.700 8.700 154.800 ;
        RECT 7.500 154.200 7.900 154.300 ;
        RECT 11.700 154.200 12.000 156.100 ;
        RECT 14.300 155.800 14.600 157.500 ;
        RECT 16.900 156.400 17.300 159.900 ;
        RECT 19.000 157.500 19.400 159.500 ;
        RECT 21.700 159.200 22.100 159.900 ;
        RECT 21.400 158.800 22.100 159.200 ;
        RECT 12.700 155.500 14.600 155.800 ;
        RECT 16.500 156.100 17.300 156.400 ;
        RECT 12.700 154.500 13.000 155.500 ;
        RECT 3.900 153.900 9.400 154.200 ;
        RECT 4.100 153.800 4.500 153.900 ;
        RECT 0.600 153.300 2.500 153.600 ;
        RECT 0.600 151.100 1.000 153.300 ;
        RECT 2.100 153.200 2.500 153.300 ;
        RECT 7.000 153.200 7.300 153.900 ;
        RECT 8.600 153.800 9.400 153.900 ;
        RECT 11.000 153.800 12.000 154.200 ;
        RECT 12.300 154.100 13.000 154.500 ;
        RECT 13.400 154.400 13.800 155.200 ;
        RECT 14.200 154.400 14.600 155.200 ;
        RECT 15.800 154.800 16.200 155.600 ;
        RECT 16.500 154.200 16.800 156.100 ;
        RECT 19.100 155.800 19.400 157.500 ;
        RECT 21.700 156.400 22.100 158.800 ;
        RECT 23.800 157.500 24.200 159.500 ;
        RECT 26.500 159.200 26.900 159.900 ;
        RECT 26.200 158.800 26.900 159.200 ;
        RECT 17.500 155.500 19.400 155.800 ;
        RECT 21.300 156.100 22.100 156.400 ;
        RECT 17.500 154.500 17.800 155.500 ;
        RECT 11.700 153.500 12.000 153.800 ;
        RECT 12.500 153.900 13.000 154.100 ;
        RECT 15.000 154.100 15.400 154.200 ;
        RECT 15.800 154.100 16.800 154.200 ;
        RECT 17.100 154.100 17.800 154.500 ;
        RECT 18.200 154.400 18.600 155.200 ;
        RECT 19.000 154.400 19.400 155.200 ;
        RECT 20.600 154.800 21.000 155.600 ;
        RECT 21.300 154.200 21.600 156.100 ;
        RECT 23.900 155.800 24.200 157.500 ;
        RECT 26.500 156.400 26.900 158.800 ;
        RECT 28.600 157.500 29.000 159.500 ;
        RECT 22.300 155.500 24.200 155.800 ;
        RECT 26.100 156.100 26.900 156.400 ;
        RECT 22.300 154.500 22.600 155.500 ;
        RECT 12.500 153.600 14.600 153.900 ;
        RECT 15.000 153.800 16.800 154.100 ;
        RECT 6.100 152.700 6.500 152.800 ;
        RECT 3.000 152.100 3.400 152.500 ;
        RECT 5.100 152.400 6.500 152.700 ;
        RECT 7.000 152.400 7.400 153.200 ;
        RECT 5.100 152.100 5.400 152.400 ;
        RECT 7.800 152.100 8.200 152.500 ;
        RECT 2.700 151.800 3.400 152.100 ;
        RECT 2.700 151.100 3.300 151.800 ;
        RECT 5.000 151.100 5.400 152.100 ;
        RECT 7.200 151.800 8.200 152.100 ;
        RECT 7.200 151.100 7.600 151.800 ;
        RECT 9.400 151.100 9.800 153.500 ;
        RECT 11.700 153.300 12.100 153.500 ;
        RECT 11.700 153.000 12.500 153.300 ;
        RECT 12.100 151.500 12.500 153.000 ;
        RECT 14.300 152.500 14.600 153.600 ;
        RECT 16.500 153.500 16.800 153.800 ;
        RECT 17.300 153.900 17.800 154.100 ;
        RECT 17.300 153.600 19.400 153.900 ;
        RECT 20.600 153.800 21.600 154.200 ;
        RECT 21.900 154.100 22.600 154.500 ;
        RECT 23.000 154.400 23.400 155.200 ;
        RECT 23.800 154.400 24.200 155.200 ;
        RECT 25.400 154.800 25.800 155.600 ;
        RECT 26.100 154.200 26.400 156.100 ;
        RECT 28.700 155.800 29.000 157.500 ;
        RECT 27.100 155.500 29.000 155.800 ;
        RECT 29.400 155.600 29.800 159.900 ;
        RECT 31.500 157.900 32.100 159.900 ;
        RECT 33.800 157.900 34.200 159.900 ;
        RECT 36.000 158.200 36.400 159.900 ;
        RECT 36.000 157.900 37.000 158.200 ;
        RECT 31.800 157.500 32.200 157.900 ;
        RECT 33.900 157.600 34.200 157.900 ;
        RECT 33.500 157.300 35.300 157.600 ;
        RECT 36.600 157.500 37.000 157.900 ;
        RECT 33.500 157.200 33.900 157.300 ;
        RECT 34.900 157.200 35.300 157.300 ;
        RECT 31.000 157.000 31.700 157.200 ;
        RECT 31.000 156.800 32.100 157.000 ;
        RECT 31.400 156.600 32.100 156.800 ;
        RECT 31.800 156.100 32.100 156.600 ;
        RECT 32.900 156.500 34.000 156.800 ;
        RECT 32.900 156.400 33.300 156.500 ;
        RECT 31.800 155.800 33.000 156.100 ;
        RECT 27.100 154.500 27.400 155.500 ;
        RECT 29.400 155.300 31.500 155.600 ;
        RECT 16.500 153.300 16.900 153.500 ;
        RECT 16.500 153.000 17.300 153.300 ;
        RECT 14.200 151.500 14.600 152.500 ;
        RECT 16.900 151.500 17.300 153.000 ;
        RECT 19.100 152.500 19.400 153.600 ;
        RECT 21.300 153.500 21.600 153.800 ;
        RECT 22.100 153.900 22.600 154.100 ;
        RECT 22.100 153.600 24.200 153.900 ;
        RECT 25.400 153.800 26.400 154.200 ;
        RECT 26.700 154.100 27.400 154.500 ;
        RECT 27.800 154.400 28.200 155.200 ;
        RECT 28.600 154.400 29.000 155.200 ;
        RECT 21.300 153.300 21.700 153.500 ;
        RECT 21.300 153.000 22.100 153.300 ;
        RECT 19.000 151.500 19.400 152.500 ;
        RECT 21.700 151.500 22.100 153.000 ;
        RECT 23.900 152.500 24.200 153.600 ;
        RECT 26.100 153.500 26.400 153.800 ;
        RECT 26.900 153.900 27.400 154.100 ;
        RECT 26.900 153.600 29.000 153.900 ;
        RECT 26.100 153.300 26.500 153.500 ;
        RECT 26.100 153.000 26.900 153.300 ;
        RECT 23.800 151.500 24.200 152.500 ;
        RECT 26.500 151.500 26.900 153.000 ;
        RECT 28.700 152.500 29.000 153.600 ;
        RECT 28.600 151.500 29.000 152.500 ;
        RECT 29.400 153.600 29.800 155.300 ;
        RECT 31.100 155.200 31.500 155.300 ;
        RECT 30.300 154.900 30.700 155.000 ;
        RECT 30.300 154.600 32.200 154.900 ;
        RECT 31.800 154.500 32.200 154.600 ;
        RECT 32.700 154.200 33.000 155.800 ;
        RECT 33.700 155.900 34.000 156.500 ;
        RECT 34.300 156.500 34.700 156.600 ;
        RECT 36.600 156.500 37.000 156.600 ;
        RECT 34.300 156.200 37.000 156.500 ;
        RECT 33.700 155.700 36.100 155.900 ;
        RECT 38.200 155.700 38.600 159.900 ;
        RECT 33.700 155.600 38.600 155.700 ;
        RECT 35.700 155.500 38.600 155.600 ;
        RECT 35.800 155.400 38.600 155.500 ;
        RECT 39.000 155.700 39.400 159.900 ;
        RECT 41.200 158.200 41.600 159.900 ;
        RECT 40.600 157.900 41.600 158.200 ;
        RECT 43.400 157.900 43.800 159.900 ;
        RECT 45.500 157.900 46.100 159.900 ;
        RECT 40.600 157.500 41.000 157.900 ;
        RECT 43.400 157.600 43.700 157.900 ;
        RECT 42.300 157.300 44.100 157.600 ;
        RECT 45.400 157.500 45.800 157.900 ;
        RECT 42.300 157.200 42.700 157.300 ;
        RECT 43.700 157.200 44.100 157.300 ;
        RECT 40.600 156.500 41.000 156.600 ;
        RECT 42.900 156.500 43.300 156.600 ;
        RECT 40.600 156.200 43.300 156.500 ;
        RECT 43.600 156.500 44.700 156.800 ;
        RECT 43.600 155.900 43.900 156.500 ;
        RECT 44.300 156.400 44.700 156.500 ;
        RECT 45.500 156.600 46.200 157.000 ;
        RECT 45.500 156.100 45.800 156.600 ;
        RECT 41.500 155.700 43.900 155.900 ;
        RECT 39.000 155.600 43.900 155.700 ;
        RECT 44.600 155.800 45.800 156.100 ;
        RECT 39.000 155.500 41.900 155.600 ;
        RECT 39.000 155.400 41.800 155.500 ;
        RECT 35.000 155.100 35.400 155.200 ;
        RECT 42.200 155.100 42.600 155.200 ;
        RECT 35.000 154.800 37.500 155.100 ;
        RECT 35.800 154.700 36.200 154.800 ;
        RECT 37.100 154.700 37.500 154.800 ;
        RECT 40.100 154.800 42.600 155.100 ;
        RECT 40.100 154.700 40.500 154.800 ;
        RECT 41.400 154.700 41.800 154.800 ;
        RECT 36.300 154.200 36.700 154.300 ;
        RECT 40.900 154.200 41.300 154.300 ;
        RECT 44.600 154.200 44.900 155.800 ;
        RECT 47.800 155.600 48.200 159.900 ;
        RECT 46.100 155.300 48.200 155.600 ;
        RECT 46.100 155.200 46.500 155.300 ;
        RECT 46.900 154.900 47.300 155.000 ;
        RECT 45.400 154.600 47.300 154.900 ;
        RECT 45.400 154.500 45.800 154.600 ;
        RECT 32.600 153.900 38.200 154.200 ;
        RECT 32.600 153.800 33.300 153.900 ;
        RECT 29.400 153.300 31.300 153.600 ;
        RECT 29.400 151.100 29.800 153.300 ;
        RECT 30.900 153.200 31.300 153.300 ;
        RECT 35.800 152.800 36.100 153.900 ;
        RECT 37.400 153.800 38.200 153.900 ;
        RECT 39.400 153.900 44.900 154.200 ;
        RECT 39.400 153.800 40.200 153.900 ;
        RECT 34.900 152.700 35.300 152.800 ;
        RECT 31.800 152.100 32.200 152.500 ;
        RECT 33.900 152.400 35.300 152.700 ;
        RECT 35.800 152.400 36.200 152.800 ;
        RECT 33.900 152.100 34.200 152.400 ;
        RECT 36.600 152.100 37.000 152.500 ;
        RECT 31.500 151.800 32.200 152.100 ;
        RECT 31.500 151.100 32.100 151.800 ;
        RECT 33.800 151.100 34.200 152.100 ;
        RECT 36.000 151.800 37.000 152.100 ;
        RECT 36.000 151.100 36.400 151.800 ;
        RECT 38.200 151.100 38.600 153.500 ;
        RECT 39.000 151.100 39.400 153.500 ;
        RECT 41.500 152.800 41.800 153.900 ;
        RECT 42.200 153.800 42.600 153.900 ;
        RECT 44.300 153.800 44.700 153.900 ;
        RECT 47.800 153.600 48.200 155.300 ;
        RECT 46.300 153.300 48.200 153.600 ;
        RECT 46.300 153.200 46.700 153.300 ;
        RECT 40.600 152.100 41.000 152.500 ;
        RECT 41.400 152.400 41.800 152.800 ;
        RECT 42.300 152.700 42.700 152.800 ;
        RECT 42.300 152.400 43.700 152.700 ;
        RECT 43.400 152.100 43.700 152.400 ;
        RECT 45.400 152.100 45.800 152.500 ;
        RECT 40.600 151.800 41.600 152.100 ;
        RECT 41.200 151.100 41.600 151.800 ;
        RECT 43.400 151.100 43.800 152.100 ;
        RECT 45.400 151.800 46.100 152.100 ;
        RECT 45.500 151.100 46.100 151.800 ;
        RECT 47.800 151.100 48.200 153.300 ;
        RECT 50.200 151.100 50.600 159.900 ;
        RECT 51.800 155.600 52.200 159.900 ;
        RECT 53.900 157.900 54.500 159.900 ;
        RECT 56.200 157.900 56.600 159.900 ;
        RECT 58.400 158.200 58.800 159.900 ;
        RECT 58.400 157.900 59.400 158.200 ;
        RECT 54.200 157.500 54.600 157.900 ;
        RECT 56.300 157.600 56.600 157.900 ;
        RECT 55.900 157.300 57.700 157.600 ;
        RECT 59.000 157.500 59.400 157.900 ;
        RECT 55.900 157.200 56.300 157.300 ;
        RECT 57.300 157.200 57.700 157.300 ;
        RECT 53.800 156.600 54.500 157.000 ;
        RECT 54.200 156.100 54.500 156.600 ;
        RECT 55.300 156.500 56.400 156.800 ;
        RECT 55.300 156.400 55.700 156.500 ;
        RECT 54.200 155.800 55.400 156.100 ;
        RECT 51.800 155.300 53.900 155.600 ;
        RECT 51.800 153.600 52.200 155.300 ;
        RECT 53.500 155.200 53.900 155.300 ;
        RECT 55.100 155.200 55.400 155.800 ;
        RECT 56.100 155.900 56.400 156.500 ;
        RECT 56.700 156.500 57.100 156.600 ;
        RECT 59.000 156.500 59.400 156.600 ;
        RECT 56.700 156.200 59.400 156.500 ;
        RECT 56.100 155.700 58.500 155.900 ;
        RECT 60.600 155.700 61.000 159.900 ;
        RECT 56.100 155.600 61.000 155.700 ;
        RECT 58.100 155.500 61.000 155.600 ;
        RECT 58.200 155.400 61.000 155.500 ;
        RECT 61.400 155.600 61.800 159.900 ;
        RECT 63.500 157.900 64.100 159.900 ;
        RECT 65.800 157.900 66.200 159.900 ;
        RECT 68.000 158.200 68.400 159.900 ;
        RECT 68.000 157.900 69.000 158.200 ;
        RECT 63.800 157.500 64.200 157.900 ;
        RECT 65.900 157.600 66.200 157.900 ;
        RECT 65.500 157.300 67.300 157.600 ;
        RECT 68.600 157.500 69.000 157.900 ;
        RECT 65.500 157.200 65.900 157.300 ;
        RECT 66.900 157.200 67.300 157.300 ;
        RECT 63.400 156.600 64.100 157.000 ;
        RECT 63.800 156.100 64.100 156.600 ;
        RECT 64.900 156.500 66.000 156.800 ;
        RECT 64.900 156.400 65.300 156.500 ;
        RECT 63.800 155.800 65.000 156.100 ;
        RECT 61.400 155.300 63.500 155.600 ;
        RECT 52.700 154.900 53.100 155.000 ;
        RECT 52.700 154.600 54.600 154.900 ;
        RECT 55.000 154.800 55.400 155.200 ;
        RECT 57.400 155.100 57.800 155.200 ;
        RECT 57.400 154.800 59.900 155.100 ;
        RECT 54.200 154.500 54.600 154.600 ;
        RECT 55.100 154.200 55.400 154.800 ;
        RECT 59.500 154.700 59.900 154.800 ;
        RECT 58.700 154.200 59.100 154.300 ;
        RECT 55.100 153.900 60.600 154.200 ;
        RECT 55.300 153.800 55.700 153.900 ;
        RECT 51.800 153.300 53.700 153.600 ;
        RECT 51.000 152.400 51.400 153.200 ;
        RECT 51.800 151.100 52.200 153.300 ;
        RECT 53.300 153.200 53.700 153.300 ;
        RECT 58.200 152.800 58.500 153.900 ;
        RECT 59.800 153.800 60.600 153.900 ;
        RECT 61.400 153.600 61.800 155.300 ;
        RECT 63.100 155.200 63.500 155.300 ;
        RECT 62.300 154.900 62.700 155.000 ;
        RECT 62.300 154.600 64.200 154.900 ;
        RECT 63.800 154.500 64.200 154.600 ;
        RECT 64.700 154.200 65.000 155.800 ;
        RECT 65.700 155.900 66.000 156.500 ;
        RECT 66.300 156.500 66.700 156.600 ;
        RECT 68.600 156.500 69.000 156.600 ;
        RECT 66.300 156.200 69.000 156.500 ;
        RECT 65.700 155.700 68.100 155.900 ;
        RECT 70.200 155.700 70.600 159.900 ;
        RECT 65.700 155.600 70.600 155.700 ;
        RECT 67.700 155.500 70.600 155.600 ;
        RECT 67.800 155.400 70.600 155.500 ;
        RECT 71.000 155.600 71.400 159.900 ;
        RECT 73.100 157.900 73.700 159.900 ;
        RECT 75.400 157.900 75.800 159.900 ;
        RECT 77.600 158.200 78.000 159.900 ;
        RECT 77.600 157.900 78.600 158.200 ;
        RECT 73.400 157.500 73.800 157.900 ;
        RECT 75.500 157.600 75.800 157.900 ;
        RECT 75.100 157.300 76.900 157.600 ;
        RECT 78.200 157.500 78.600 157.900 ;
        RECT 75.100 157.200 75.500 157.300 ;
        RECT 76.500 157.200 76.900 157.300 ;
        RECT 73.000 156.600 73.700 157.000 ;
        RECT 73.400 156.100 73.700 156.600 ;
        RECT 74.500 156.500 75.600 156.800 ;
        RECT 74.500 156.400 74.900 156.500 ;
        RECT 73.400 155.800 74.600 156.100 ;
        RECT 71.000 155.300 73.100 155.600 ;
        RECT 67.000 155.100 67.400 155.200 ;
        RECT 67.000 154.800 69.500 155.100 ;
        RECT 69.100 154.700 69.500 154.800 ;
        RECT 68.300 154.200 68.700 154.300 ;
        RECT 64.700 153.900 70.200 154.200 ;
        RECT 64.900 153.800 65.300 153.900 ;
        RECT 57.300 152.700 57.700 152.800 ;
        RECT 54.200 152.100 54.600 152.500 ;
        RECT 56.300 152.400 57.700 152.700 ;
        RECT 58.200 152.400 58.600 152.800 ;
        RECT 56.300 152.100 56.600 152.400 ;
        RECT 59.000 152.100 59.400 152.500 ;
        RECT 53.900 151.800 54.600 152.100 ;
        RECT 53.900 151.100 54.500 151.800 ;
        RECT 56.200 151.100 56.600 152.100 ;
        RECT 58.400 151.800 59.400 152.100 ;
        RECT 58.400 151.100 58.800 151.800 ;
        RECT 60.600 151.100 61.000 153.500 ;
        RECT 61.400 153.300 63.300 153.600 ;
        RECT 61.400 151.100 61.800 153.300 ;
        RECT 62.900 153.200 63.300 153.300 ;
        RECT 67.800 152.800 68.100 153.900 ;
        RECT 69.400 153.800 70.200 153.900 ;
        RECT 71.000 153.600 71.400 155.300 ;
        RECT 72.700 155.200 73.100 155.300 ;
        RECT 71.900 154.900 72.300 155.000 ;
        RECT 71.900 154.600 73.800 154.900 ;
        RECT 73.400 154.500 73.800 154.600 ;
        RECT 74.300 154.200 74.600 155.800 ;
        RECT 75.300 155.900 75.600 156.500 ;
        RECT 75.900 156.500 76.300 156.600 ;
        RECT 78.200 156.500 78.600 156.600 ;
        RECT 75.900 156.200 78.600 156.500 ;
        RECT 75.300 155.700 77.700 155.900 ;
        RECT 79.800 155.700 80.200 159.900 ;
        RECT 75.300 155.600 80.200 155.700 ;
        RECT 77.300 155.500 80.200 155.600 ;
        RECT 77.400 155.400 80.200 155.500 ;
        RECT 80.600 155.600 81.000 159.900 ;
        RECT 82.700 157.900 83.300 159.900 ;
        RECT 85.000 157.900 85.400 159.900 ;
        RECT 87.200 158.200 87.600 159.900 ;
        RECT 87.200 157.900 88.200 158.200 ;
        RECT 83.000 157.500 83.400 157.900 ;
        RECT 85.100 157.600 85.400 157.900 ;
        RECT 84.700 157.300 86.500 157.600 ;
        RECT 87.800 157.500 88.200 157.900 ;
        RECT 84.700 157.200 85.100 157.300 ;
        RECT 86.100 157.200 86.500 157.300 ;
        RECT 82.200 157.000 82.900 157.200 ;
        RECT 82.200 156.800 83.300 157.000 ;
        RECT 82.600 156.600 83.300 156.800 ;
        RECT 83.000 156.100 83.300 156.600 ;
        RECT 84.100 156.500 85.200 156.800 ;
        RECT 84.100 156.400 84.500 156.500 ;
        RECT 83.000 155.800 84.200 156.100 ;
        RECT 80.600 155.300 82.700 155.600 ;
        RECT 76.600 155.100 77.000 155.200 ;
        RECT 76.600 154.800 79.100 155.100 ;
        RECT 77.400 154.700 77.800 154.800 ;
        RECT 78.700 154.700 79.100 154.800 ;
        RECT 77.900 154.200 78.300 154.300 ;
        RECT 74.300 153.900 79.800 154.200 ;
        RECT 74.500 153.800 74.900 153.900 ;
        RECT 66.900 152.700 67.300 152.800 ;
        RECT 63.800 152.100 64.200 152.500 ;
        RECT 65.900 152.400 67.300 152.700 ;
        RECT 67.800 152.400 68.200 152.800 ;
        RECT 65.900 152.100 66.200 152.400 ;
        RECT 68.600 152.100 69.000 152.500 ;
        RECT 63.500 151.800 64.200 152.100 ;
        RECT 63.500 151.100 64.100 151.800 ;
        RECT 65.800 151.100 66.200 152.100 ;
        RECT 68.000 151.800 69.000 152.100 ;
        RECT 68.000 151.100 68.400 151.800 ;
        RECT 70.200 151.100 70.600 153.500 ;
        RECT 71.000 153.300 72.900 153.600 ;
        RECT 71.000 151.100 71.400 153.300 ;
        RECT 72.500 153.200 72.900 153.300 ;
        RECT 77.400 153.200 77.700 153.900 ;
        RECT 79.000 153.800 79.800 153.900 ;
        RECT 80.600 153.600 81.000 155.300 ;
        RECT 82.300 155.200 82.700 155.300 ;
        RECT 81.500 154.900 81.900 155.000 ;
        RECT 81.500 154.600 83.400 154.900 ;
        RECT 83.000 154.500 83.400 154.600 ;
        RECT 83.900 154.200 84.200 155.800 ;
        RECT 84.900 155.900 85.200 156.500 ;
        RECT 85.500 156.500 85.900 156.600 ;
        RECT 87.800 156.500 88.200 156.600 ;
        RECT 85.500 156.200 88.200 156.500 ;
        RECT 84.900 155.700 87.300 155.900 ;
        RECT 89.400 155.700 89.800 159.900 ;
        RECT 92.100 156.400 92.500 159.900 ;
        RECT 94.200 157.500 94.600 159.500 ;
        RECT 84.900 155.600 89.800 155.700 ;
        RECT 91.700 156.100 92.500 156.400 ;
        RECT 86.900 155.500 89.800 155.600 ;
        RECT 87.000 155.400 89.800 155.500 ;
        RECT 86.200 155.100 86.600 155.200 ;
        RECT 86.200 154.800 88.700 155.100 ;
        RECT 91.000 154.800 91.400 155.600 ;
        RECT 87.000 154.700 87.400 154.800 ;
        RECT 88.300 154.700 88.700 154.800 ;
        RECT 87.500 154.200 87.900 154.300 ;
        RECT 91.700 154.200 92.000 156.100 ;
        RECT 94.300 155.800 94.600 157.500 ;
        RECT 95.000 156.200 95.400 159.900 ;
        RECT 96.600 156.200 97.000 159.900 ;
        RECT 95.000 155.900 97.000 156.200 ;
        RECT 97.400 157.100 97.800 159.900 ;
        RECT 98.200 157.100 98.600 157.200 ;
        RECT 97.400 156.800 98.600 157.100 ;
        RECT 97.400 155.900 97.800 156.800 ;
        RECT 101.100 156.200 101.500 159.900 ;
        RECT 101.800 156.800 102.200 157.200 ;
        RECT 101.900 156.200 102.200 156.800 ;
        RECT 103.300 156.300 103.700 159.900 ;
        RECT 101.100 155.900 101.600 156.200 ;
        RECT 101.900 155.900 102.600 156.200 ;
        RECT 103.300 155.900 104.200 156.300 ;
        RECT 105.400 156.200 105.800 159.900 ;
        RECT 107.800 156.200 108.200 159.900 ;
        RECT 110.200 157.500 110.600 159.500 ;
        RECT 112.300 159.200 112.700 159.900 ;
        RECT 111.800 158.800 112.700 159.200 ;
        RECT 105.400 155.900 106.500 156.200 ;
        RECT 107.800 155.900 108.900 156.200 ;
        RECT 92.700 155.500 94.600 155.800 ;
        RECT 92.700 154.500 93.000 155.500 ;
        RECT 95.400 155.200 95.800 155.400 ;
        RECT 97.400 155.200 97.700 155.900 ;
        RECT 101.300 155.200 101.600 155.900 ;
        RECT 102.200 155.800 102.600 155.900 ;
        RECT 83.900 153.900 89.400 154.200 ;
        RECT 84.100 153.800 84.500 153.900 ;
        RECT 76.500 152.700 76.900 152.800 ;
        RECT 73.400 152.100 73.800 152.500 ;
        RECT 75.500 152.400 76.900 152.700 ;
        RECT 77.400 152.400 77.800 153.200 ;
        RECT 75.500 152.100 75.800 152.400 ;
        RECT 78.200 152.100 78.600 152.500 ;
        RECT 73.100 151.800 73.800 152.100 ;
        RECT 73.100 151.100 73.700 151.800 ;
        RECT 75.400 151.100 75.800 152.100 ;
        RECT 77.600 151.800 78.600 152.100 ;
        RECT 77.600 151.100 78.000 151.800 ;
        RECT 79.800 151.100 80.200 153.500 ;
        RECT 80.600 153.300 82.500 153.600 ;
        RECT 80.600 151.100 81.000 153.300 ;
        RECT 82.100 153.200 82.500 153.300 ;
        RECT 87.000 152.800 87.300 153.900 ;
        RECT 88.600 153.800 89.400 153.900 ;
        RECT 91.000 153.800 92.000 154.200 ;
        RECT 92.300 154.100 93.000 154.500 ;
        RECT 93.400 154.400 93.800 155.200 ;
        RECT 94.200 154.400 94.600 155.200 ;
        RECT 95.000 154.900 95.800 155.200 ;
        RECT 96.600 154.900 97.800 155.200 ;
        RECT 95.000 154.800 95.400 154.900 ;
        RECT 91.700 153.500 92.000 153.800 ;
        RECT 92.500 153.900 93.000 154.100 ;
        RECT 92.500 153.600 94.600 153.900 ;
        RECT 95.800 153.800 96.200 154.600 ;
        RECT 86.100 152.700 86.500 152.800 ;
        RECT 83.000 152.100 83.400 152.500 ;
        RECT 85.100 152.400 86.500 152.700 ;
        RECT 87.000 152.400 87.400 152.800 ;
        RECT 85.100 152.100 85.400 152.400 ;
        RECT 87.800 152.100 88.200 152.500 ;
        RECT 82.700 151.800 83.400 152.100 ;
        RECT 82.700 151.100 83.300 151.800 ;
        RECT 85.000 151.100 85.400 152.100 ;
        RECT 87.200 151.800 88.200 152.100 ;
        RECT 87.200 151.100 87.600 151.800 ;
        RECT 89.400 151.100 89.800 153.500 ;
        RECT 91.700 153.300 92.100 153.500 ;
        RECT 91.700 153.200 92.500 153.300 ;
        RECT 91.700 153.000 93.000 153.200 ;
        RECT 92.100 152.800 93.000 153.000 ;
        RECT 92.100 151.500 92.500 152.800 ;
        RECT 94.300 152.500 94.600 153.600 ;
        RECT 94.200 151.500 94.600 152.500 ;
        RECT 96.600 153.100 96.900 154.900 ;
        RECT 97.400 154.800 97.800 154.900 ;
        RECT 100.600 154.400 101.000 155.200 ;
        RECT 101.300 154.800 101.800 155.200 ;
        RECT 103.000 154.800 103.400 155.600 ;
        RECT 103.800 155.100 104.100 155.900 ;
        RECT 106.200 155.600 106.500 155.900 ;
        RECT 108.600 155.600 108.900 155.900 ;
        RECT 110.200 155.800 110.500 157.500 ;
        RECT 112.300 156.400 112.700 158.800 ;
        RECT 112.300 156.100 113.100 156.400 ;
        RECT 116.600 156.200 117.000 159.900 ;
        RECT 118.700 156.300 119.100 159.900 ;
        RECT 106.200 155.200 106.800 155.600 ;
        RECT 108.600 155.200 109.200 155.600 ;
        RECT 110.200 155.500 112.100 155.800 ;
        RECT 105.400 155.100 105.800 155.200 ;
        RECT 103.800 154.800 105.800 155.100 ;
        RECT 101.300 154.200 101.600 154.800 ;
        RECT 103.800 154.200 104.100 154.800 ;
        RECT 105.400 154.400 105.800 154.800 ;
        RECT 99.800 154.100 100.200 154.200 ;
        RECT 97.400 153.800 100.600 154.100 ;
        RECT 101.300 153.800 102.600 154.200 ;
        RECT 103.800 153.800 104.200 154.200 ;
        RECT 97.400 153.200 97.700 153.800 ;
        RECT 100.200 153.600 100.600 153.800 ;
        RECT 96.600 151.100 97.000 153.100 ;
        RECT 97.400 152.800 97.800 153.200 ;
        RECT 99.900 153.100 101.700 153.300 ;
        RECT 102.200 153.100 102.500 153.800 ;
        RECT 99.800 153.000 101.800 153.100 ;
        RECT 97.300 152.400 97.700 152.800 ;
        RECT 99.800 151.100 100.200 153.000 ;
        RECT 101.400 151.100 101.800 153.000 ;
        RECT 102.200 151.100 102.600 153.100 ;
        RECT 103.800 152.100 104.100 153.800 ;
        RECT 106.200 153.700 106.500 155.200 ;
        RECT 107.800 154.400 108.200 155.200 ;
        RECT 108.600 153.700 108.900 155.200 ;
        RECT 110.200 154.400 110.600 155.200 ;
        RECT 111.000 154.400 111.400 155.200 ;
        RECT 111.800 154.500 112.100 155.500 ;
        RECT 111.800 154.100 112.500 154.500 ;
        RECT 112.800 154.200 113.100 156.100 ;
        RECT 115.900 155.900 117.000 156.200 ;
        RECT 118.200 155.900 119.100 156.300 ;
        RECT 119.800 155.900 120.200 159.900 ;
        RECT 120.600 156.200 121.000 159.900 ;
        RECT 122.200 156.200 122.600 159.900 ;
        RECT 123.400 156.800 123.800 157.200 ;
        RECT 123.400 156.200 123.700 156.800 ;
        RECT 124.100 156.200 124.500 159.900 ;
        RECT 120.600 155.900 122.600 156.200 ;
        RECT 123.000 155.900 123.700 156.200 ;
        RECT 124.000 155.900 124.500 156.200 ;
        RECT 115.900 155.600 116.200 155.900 ;
        RECT 113.400 154.800 113.800 155.600 ;
        RECT 115.600 155.200 116.200 155.600 ;
        RECT 111.800 153.900 112.300 154.100 ;
        RECT 105.400 153.400 106.500 153.700 ;
        RECT 107.800 153.400 108.900 153.700 ;
        RECT 110.200 153.600 112.300 153.900 ;
        RECT 112.800 153.800 113.800 154.200 ;
        RECT 104.600 152.400 105.000 153.200 ;
        RECT 103.800 151.100 104.200 152.100 ;
        RECT 105.400 151.100 105.800 153.400 ;
        RECT 107.800 151.100 108.200 153.400 ;
        RECT 110.200 152.500 110.500 153.600 ;
        RECT 112.800 153.500 113.100 153.800 ;
        RECT 112.700 153.300 113.100 153.500 ;
        RECT 115.900 153.700 116.200 155.200 ;
        RECT 116.600 155.100 117.000 155.200 ;
        RECT 118.300 155.100 118.600 155.900 ;
        RECT 116.600 154.800 118.600 155.100 ;
        RECT 119.000 155.100 119.400 155.600 ;
        RECT 119.900 155.200 120.200 155.900 ;
        RECT 123.000 155.800 123.400 155.900 ;
        RECT 121.800 155.200 122.200 155.400 ;
        RECT 119.800 155.100 121.000 155.200 ;
        RECT 119.000 154.900 121.000 155.100 ;
        RECT 121.800 155.100 122.600 155.200 ;
        RECT 123.000 155.100 123.300 155.800 ;
        RECT 124.000 155.200 124.300 155.900 ;
        RECT 121.800 154.900 123.300 155.100 ;
        RECT 119.000 154.800 120.200 154.900 ;
        RECT 116.600 154.400 117.000 154.800 ;
        RECT 118.300 154.200 118.600 154.800 ;
        RECT 118.200 153.800 118.600 154.200 ;
        RECT 115.900 153.400 117.000 153.700 ;
        RECT 112.300 153.000 113.100 153.300 ;
        RECT 110.200 151.500 110.600 152.500 ;
        RECT 112.300 151.500 112.700 153.000 ;
        RECT 116.600 151.100 117.000 153.400 ;
        RECT 117.400 152.400 117.800 153.200 ;
        RECT 118.300 152.100 118.600 153.800 ;
        RECT 119.800 152.800 120.200 153.200 ;
        RECT 120.700 153.100 121.000 154.900 ;
        RECT 122.200 154.800 123.300 154.900 ;
        RECT 123.800 154.800 124.300 155.200 ;
        RECT 121.400 153.800 121.800 154.600 ;
        RECT 124.000 154.200 124.300 154.800 ;
        RECT 124.600 155.100 125.000 155.200 ;
        RECT 125.400 155.100 125.800 155.200 ;
        RECT 124.600 154.800 125.800 155.100 ;
        RECT 124.600 154.400 125.000 154.800 ;
        RECT 123.000 153.800 124.300 154.200 ;
        RECT 125.400 154.100 125.800 154.200 ;
        RECT 125.000 153.800 126.500 154.100 ;
        RECT 123.100 153.100 123.400 153.800 ;
        RECT 125.000 153.600 125.400 153.800 ;
        RECT 123.900 153.100 125.700 153.300 ;
        RECT 126.200 153.200 126.500 153.800 ;
        RECT 119.900 152.400 120.300 152.800 ;
        RECT 118.200 151.100 118.600 152.100 ;
        RECT 120.600 151.100 121.000 153.100 ;
        RECT 123.000 151.100 123.400 153.100 ;
        RECT 123.800 153.000 125.800 153.100 ;
        RECT 123.800 151.100 124.200 153.000 ;
        RECT 125.400 151.100 125.800 153.000 ;
        RECT 126.200 152.400 126.600 153.200 ;
        RECT 127.000 151.100 127.400 159.900 ;
        RECT 129.100 156.300 129.500 159.900 ;
        RECT 128.600 155.900 129.500 156.300 ;
        RECT 130.200 156.200 130.600 159.900 ;
        RECT 132.900 156.300 133.300 159.900 ;
        RECT 130.200 155.900 131.300 156.200 ;
        RECT 132.900 155.900 133.800 156.300 ;
        RECT 128.700 155.200 129.000 155.900 ;
        RECT 131.000 155.600 131.300 155.900 ;
        RECT 128.600 154.800 129.000 155.200 ;
        RECT 129.400 154.800 129.800 155.600 ;
        RECT 131.000 155.200 131.600 155.600 ;
        RECT 128.700 154.200 129.000 154.800 ;
        RECT 130.200 154.400 130.600 155.200 ;
        RECT 128.600 153.800 129.000 154.200 ;
        RECT 127.800 152.400 128.200 153.200 ;
        RECT 128.700 152.100 129.000 153.800 ;
        RECT 131.000 153.700 131.300 155.200 ;
        RECT 132.600 154.800 133.000 155.600 ;
        RECT 133.400 155.100 133.700 155.900 ;
        RECT 135.000 155.600 135.400 159.900 ;
        RECT 137.100 157.900 137.700 159.900 ;
        RECT 139.400 157.900 139.800 159.900 ;
        RECT 141.600 158.200 142.000 159.900 ;
        RECT 141.600 157.900 142.600 158.200 ;
        RECT 137.400 157.500 137.800 157.900 ;
        RECT 139.500 157.600 139.800 157.900 ;
        RECT 139.100 157.300 140.900 157.600 ;
        RECT 142.200 157.500 142.600 157.900 ;
        RECT 139.100 157.200 139.500 157.300 ;
        RECT 140.500 157.200 140.900 157.300 ;
        RECT 137.000 156.600 137.700 157.000 ;
        RECT 137.400 156.100 137.700 156.600 ;
        RECT 138.500 156.500 139.600 156.800 ;
        RECT 138.500 156.400 138.900 156.500 ;
        RECT 137.400 155.800 138.600 156.100 ;
        RECT 135.000 155.300 137.100 155.600 ;
        RECT 133.400 154.800 134.500 155.100 ;
        RECT 128.600 151.100 129.000 152.100 ;
        RECT 130.200 153.400 131.300 153.700 ;
        RECT 133.400 154.200 133.700 154.800 ;
        RECT 134.200 154.200 134.500 154.800 ;
        RECT 133.400 153.800 133.800 154.200 ;
        RECT 134.200 153.800 134.600 154.200 ;
        RECT 130.200 151.100 130.600 153.400 ;
        RECT 133.400 152.100 133.700 153.800 ;
        RECT 135.000 153.600 135.400 155.300 ;
        RECT 136.700 155.200 137.100 155.300 ;
        RECT 138.300 155.200 138.600 155.800 ;
        RECT 139.300 155.900 139.600 156.500 ;
        RECT 139.900 156.500 140.300 156.600 ;
        RECT 142.200 156.500 142.600 156.600 ;
        RECT 139.900 156.200 142.600 156.500 ;
        RECT 139.300 155.700 141.700 155.900 ;
        RECT 143.800 155.700 144.200 159.900 ;
        RECT 146.500 156.400 146.900 159.900 ;
        RECT 148.600 157.500 149.000 159.500 ;
        RECT 139.300 155.600 144.200 155.700 ;
        RECT 146.100 156.100 146.900 156.400 ;
        RECT 141.300 155.500 144.200 155.600 ;
        RECT 141.400 155.400 144.200 155.500 ;
        RECT 135.900 154.900 136.300 155.000 ;
        RECT 135.900 154.600 137.800 154.900 ;
        RECT 138.200 154.800 138.600 155.200 ;
        RECT 140.600 155.100 141.000 155.200 ;
        RECT 140.600 154.800 143.100 155.100 ;
        RECT 137.400 154.500 137.800 154.600 ;
        RECT 138.300 154.200 138.600 154.800 ;
        RECT 142.700 154.700 143.100 154.800 ;
        RECT 144.600 154.800 145.000 155.200 ;
        RECT 145.400 154.800 145.800 155.600 ;
        RECT 146.100 155.200 146.400 156.100 ;
        RECT 148.700 155.800 149.000 157.500 ;
        RECT 151.300 156.300 151.700 159.900 ;
        RECT 151.300 155.900 152.200 156.300 ;
        RECT 147.100 155.500 149.000 155.800 ;
        RECT 146.100 154.800 146.600 155.200 ;
        RECT 141.900 154.200 142.300 154.300 ;
        RECT 138.300 154.100 143.800 154.200 ;
        RECT 144.600 154.100 144.900 154.800 ;
        RECT 146.100 154.200 146.400 154.800 ;
        RECT 147.100 154.500 147.400 155.500 ;
        RECT 138.300 153.900 144.900 154.100 ;
        RECT 138.500 153.800 138.900 153.900 ;
        RECT 135.000 153.300 136.900 153.600 ;
        RECT 134.200 152.400 134.600 153.200 ;
        RECT 133.400 151.100 133.800 152.100 ;
        RECT 135.000 151.100 135.400 153.300 ;
        RECT 136.500 153.200 136.900 153.300 ;
        RECT 141.400 152.800 141.700 153.900 ;
        RECT 143.000 153.800 144.900 153.900 ;
        RECT 145.400 153.800 146.400 154.200 ;
        RECT 146.700 154.100 147.400 154.500 ;
        RECT 147.800 154.400 148.200 155.200 ;
        RECT 148.600 155.100 149.000 155.200 ;
        RECT 150.200 155.100 150.600 155.200 ;
        RECT 148.600 154.800 150.600 155.100 ;
        RECT 151.000 154.800 151.400 155.600 ;
        RECT 148.600 154.400 149.000 154.800 ;
        RECT 146.100 153.500 146.400 153.800 ;
        RECT 146.900 153.900 147.400 154.100 ;
        RECT 151.800 154.200 152.100 155.900 ;
        RECT 153.400 155.700 153.800 159.900 ;
        RECT 155.600 158.200 156.000 159.900 ;
        RECT 155.000 157.900 156.000 158.200 ;
        RECT 157.800 157.900 158.200 159.900 ;
        RECT 159.900 157.900 160.500 159.900 ;
        RECT 155.000 157.500 155.400 157.900 ;
        RECT 157.800 157.600 158.100 157.900 ;
        RECT 156.700 157.300 158.500 157.600 ;
        RECT 159.800 157.500 160.200 157.900 ;
        RECT 156.700 157.200 157.100 157.300 ;
        RECT 158.100 157.200 158.500 157.300 ;
        RECT 160.300 157.000 161.000 157.200 ;
        RECT 159.900 156.800 161.000 157.000 ;
        RECT 155.000 156.500 155.400 156.600 ;
        RECT 157.300 156.500 157.700 156.600 ;
        RECT 155.000 156.200 157.700 156.500 ;
        RECT 158.000 156.500 159.100 156.800 ;
        RECT 158.000 155.900 158.300 156.500 ;
        RECT 158.700 156.400 159.100 156.500 ;
        RECT 159.900 156.600 160.600 156.800 ;
        RECT 159.900 156.100 160.200 156.600 ;
        RECT 155.900 155.700 158.300 155.900 ;
        RECT 153.400 155.600 158.300 155.700 ;
        RECT 159.000 155.800 160.200 156.100 ;
        RECT 153.400 155.500 156.300 155.600 ;
        RECT 153.400 155.400 156.200 155.500 ;
        RECT 156.600 155.100 157.000 155.200 ;
        RECT 154.500 154.800 157.000 155.100 ;
        RECT 154.500 154.700 154.900 154.800 ;
        RECT 155.300 154.200 155.700 154.300 ;
        RECT 159.000 154.200 159.300 155.800 ;
        RECT 162.200 155.600 162.600 159.900 ;
        RECT 160.500 155.300 162.600 155.600 ;
        RECT 160.500 155.200 160.900 155.300 ;
        RECT 161.300 154.900 161.700 155.000 ;
        RECT 159.800 154.600 161.700 154.900 ;
        RECT 159.800 154.500 160.200 154.600 ;
        RECT 146.900 153.600 149.000 153.900 ;
        RECT 140.500 152.700 140.900 152.800 ;
        RECT 137.400 152.100 137.800 152.500 ;
        RECT 139.500 152.400 140.900 152.700 ;
        RECT 141.400 152.400 141.800 152.800 ;
        RECT 139.500 152.100 139.800 152.400 ;
        RECT 142.200 152.100 142.600 152.500 ;
        RECT 137.100 151.800 137.800 152.100 ;
        RECT 137.100 151.100 137.700 151.800 ;
        RECT 139.400 151.100 139.800 152.100 ;
        RECT 141.600 151.800 142.600 152.100 ;
        RECT 141.600 151.100 142.000 151.800 ;
        RECT 143.800 151.100 144.200 153.500 ;
        RECT 146.100 153.300 146.500 153.500 ;
        RECT 146.100 153.000 146.900 153.300 ;
        RECT 146.500 151.500 146.900 153.000 ;
        RECT 148.700 152.500 149.000 153.600 ;
        RECT 151.800 153.800 152.200 154.200 ;
        RECT 153.800 153.900 159.300 154.200 ;
        RECT 153.800 153.800 154.600 153.900 ;
        RECT 151.000 153.100 151.400 153.200 ;
        RECT 151.800 153.100 152.100 153.800 ;
        RECT 151.000 152.800 152.100 153.100 ;
        RECT 148.600 151.500 149.000 152.500 ;
        RECT 151.800 152.100 152.100 152.800 ;
        RECT 152.600 152.400 153.000 153.200 ;
        RECT 151.800 151.100 152.200 152.100 ;
        RECT 153.400 151.100 153.800 153.500 ;
        RECT 155.900 152.800 156.200 153.900 ;
        RECT 158.700 153.800 159.100 153.900 ;
        RECT 162.200 153.600 162.600 155.300 ;
        RECT 160.600 153.300 162.600 153.600 ;
        RECT 160.600 153.200 161.100 153.300 ;
        RECT 160.600 152.800 161.000 153.200 ;
        RECT 155.000 152.100 155.400 152.500 ;
        RECT 155.800 152.400 156.200 152.800 ;
        RECT 156.700 152.700 157.100 152.800 ;
        RECT 156.700 152.400 158.100 152.700 ;
        RECT 157.800 152.100 158.100 152.400 ;
        RECT 159.800 152.100 160.200 152.500 ;
        RECT 155.000 151.800 156.000 152.100 ;
        RECT 155.600 151.100 156.000 151.800 ;
        RECT 157.800 151.100 158.200 152.100 ;
        RECT 159.800 151.800 160.500 152.100 ;
        RECT 159.900 151.100 160.500 151.800 ;
        RECT 162.200 151.100 162.600 153.300 ;
        RECT 163.000 155.900 163.400 159.900 ;
        RECT 164.600 157.900 165.000 159.900 ;
        RECT 167.500 159.200 167.900 159.900 ;
        RECT 167.000 158.800 167.900 159.200 ;
        RECT 163.000 155.200 163.300 155.900 ;
        RECT 164.600 155.800 164.900 157.900 ;
        RECT 167.500 156.300 167.900 158.800 ;
        RECT 170.500 156.400 170.900 159.900 ;
        RECT 172.600 157.500 173.000 159.500 ;
        RECT 167.000 155.900 167.900 156.300 ;
        RECT 170.100 156.100 170.900 156.400 ;
        RECT 163.700 155.500 164.900 155.800 ;
        RECT 163.000 154.800 163.400 155.200 ;
        RECT 163.000 153.100 163.300 154.800 ;
        RECT 163.700 153.800 164.000 155.500 ;
        RECT 167.100 154.200 167.400 155.900 ;
        RECT 167.000 153.800 167.400 154.200 ;
        RECT 167.800 154.800 168.200 155.600 ;
        RECT 167.800 154.100 168.100 154.800 ;
        RECT 170.100 154.200 170.400 156.100 ;
        RECT 172.700 155.800 173.000 157.500 ;
        RECT 171.100 155.500 173.000 155.800 ;
        RECT 173.400 157.500 173.800 159.500 ;
        RECT 173.400 155.800 173.700 157.500 ;
        RECT 175.500 156.400 175.900 159.900 ;
        RECT 175.500 156.100 176.300 156.400 ;
        RECT 173.400 155.500 175.300 155.800 ;
        RECT 171.100 154.500 171.400 155.500 ;
        RECT 169.400 154.100 170.400 154.200 ;
        RECT 170.700 154.100 171.400 154.500 ;
        RECT 171.800 154.400 172.200 155.200 ;
        RECT 172.600 155.100 173.000 155.200 ;
        RECT 173.400 155.100 173.800 155.200 ;
        RECT 172.600 154.800 173.800 155.100 ;
        RECT 172.600 154.400 173.000 154.800 ;
        RECT 173.400 154.400 173.800 154.800 ;
        RECT 174.200 154.400 174.600 155.200 ;
        RECT 175.000 154.500 175.300 155.500 ;
        RECT 167.800 153.800 170.400 154.100 ;
        RECT 163.600 153.700 164.000 153.800 ;
        RECT 163.600 153.500 165.100 153.700 ;
        RECT 163.600 153.400 165.700 153.500 ;
        RECT 164.800 153.200 165.700 153.400 ;
        RECT 165.400 153.100 165.700 153.200 ;
        RECT 163.000 152.600 163.700 153.100 ;
        RECT 163.300 152.200 163.700 152.600 ;
        RECT 163.000 151.800 163.700 152.200 ;
        RECT 163.300 151.100 163.700 151.800 ;
        RECT 165.400 151.100 165.800 153.100 ;
        RECT 166.200 152.400 166.600 153.200 ;
        RECT 167.100 152.100 167.400 153.800 ;
        RECT 170.100 153.500 170.400 153.800 ;
        RECT 170.900 153.900 171.400 154.100 ;
        RECT 175.000 154.100 175.700 154.500 ;
        RECT 176.000 154.200 176.300 156.100 ;
        RECT 178.200 155.900 178.600 159.900 ;
        RECT 179.800 156.200 180.200 159.900 ;
        RECT 179.100 155.900 180.200 156.200 ;
        RECT 180.900 159.200 181.300 159.900 ;
        RECT 180.900 158.800 181.800 159.200 ;
        RECT 180.900 156.300 181.300 158.800 ;
        RECT 180.900 155.900 181.800 156.300 ;
        RECT 177.400 154.800 177.800 155.200 ;
        RECT 178.200 154.800 178.500 155.900 ;
        RECT 179.100 155.600 179.400 155.900 ;
        RECT 178.800 155.200 179.400 155.600 ;
        RECT 176.000 154.100 177.000 154.200 ;
        RECT 177.400 154.100 177.700 154.800 ;
        RECT 175.000 153.900 175.500 154.100 ;
        RECT 170.900 153.600 173.000 153.900 ;
        RECT 170.100 153.300 170.500 153.500 ;
        RECT 170.100 153.000 170.900 153.300 ;
        RECT 167.000 151.100 167.400 152.100 ;
        RECT 170.500 151.500 170.900 153.000 ;
        RECT 172.700 152.500 173.000 153.600 ;
        RECT 172.600 151.500 173.000 152.500 ;
        RECT 173.400 153.600 175.500 153.900 ;
        RECT 176.000 153.800 177.700 154.100 ;
        RECT 173.400 152.500 173.700 153.600 ;
        RECT 176.000 153.500 176.300 153.800 ;
        RECT 175.900 153.300 176.300 153.500 ;
        RECT 175.500 153.000 176.300 153.300 ;
        RECT 173.400 151.500 173.800 152.500 ;
        RECT 175.500 151.500 175.900 153.000 ;
        RECT 178.200 151.100 178.600 154.800 ;
        RECT 179.100 153.700 179.400 155.200 ;
        RECT 180.600 154.800 181.000 155.600 ;
        RECT 181.400 154.200 181.700 155.900 ;
        RECT 183.000 155.700 183.400 159.900 ;
        RECT 185.200 158.200 185.600 159.900 ;
        RECT 184.600 157.900 185.600 158.200 ;
        RECT 187.400 157.900 187.800 159.900 ;
        RECT 189.500 157.900 190.100 159.900 ;
        RECT 184.600 157.500 185.000 157.900 ;
        RECT 187.400 157.600 187.700 157.900 ;
        RECT 186.300 157.300 188.100 157.600 ;
        RECT 189.400 157.500 189.800 157.900 ;
        RECT 186.300 157.200 186.700 157.300 ;
        RECT 187.700 157.200 188.100 157.300 ;
        RECT 184.600 156.500 185.000 156.600 ;
        RECT 186.900 156.500 187.300 156.600 ;
        RECT 184.600 156.200 187.300 156.500 ;
        RECT 187.600 156.500 188.700 156.800 ;
        RECT 187.600 155.900 187.900 156.500 ;
        RECT 188.300 156.400 188.700 156.500 ;
        RECT 189.500 156.600 190.200 157.000 ;
        RECT 189.500 156.100 189.800 156.600 ;
        RECT 185.500 155.700 187.900 155.900 ;
        RECT 183.000 155.600 187.900 155.700 ;
        RECT 188.600 155.800 189.800 156.100 ;
        RECT 183.000 155.500 185.900 155.600 ;
        RECT 183.000 155.400 185.800 155.500 ;
        RECT 186.200 155.100 186.600 155.200 ;
        RECT 184.100 154.800 186.600 155.100 ;
        RECT 184.100 154.700 184.500 154.800 ;
        RECT 185.400 154.700 185.800 154.800 ;
        RECT 184.900 154.200 185.300 154.300 ;
        RECT 188.600 154.200 188.900 155.800 ;
        RECT 191.800 155.600 192.200 159.900 ;
        RECT 192.600 156.200 193.000 159.900 ;
        RECT 192.600 155.900 193.700 156.200 ;
        RECT 190.100 155.300 192.200 155.600 ;
        RECT 190.100 155.200 190.500 155.300 ;
        RECT 190.900 154.900 191.300 155.000 ;
        RECT 189.400 154.600 191.300 154.900 ;
        RECT 189.400 154.500 189.800 154.600 ;
        RECT 181.400 153.800 181.800 154.200 ;
        RECT 183.400 154.100 188.900 154.200 ;
        RECT 182.200 153.900 188.900 154.100 ;
        RECT 182.200 153.800 184.200 153.900 ;
        RECT 179.100 153.400 180.200 153.700 ;
        RECT 179.800 151.100 180.200 153.400 ;
        RECT 181.400 152.100 181.700 153.800 ;
        RECT 182.200 153.200 182.500 153.800 ;
        RECT 182.200 152.400 182.600 153.200 ;
        RECT 181.400 151.100 181.800 152.100 ;
        RECT 183.000 151.100 183.400 153.500 ;
        RECT 185.500 152.800 185.800 153.900 ;
        RECT 188.300 153.800 188.700 153.900 ;
        RECT 191.800 153.600 192.200 155.300 ;
        RECT 193.400 155.600 193.700 155.900 ;
        RECT 193.400 155.200 194.000 155.600 ;
        RECT 193.400 153.700 193.700 155.200 ;
        RECT 190.300 153.300 192.200 153.600 ;
        RECT 190.300 153.200 190.700 153.300 ;
        RECT 184.600 152.100 185.000 152.500 ;
        RECT 185.400 152.400 185.800 152.800 ;
        RECT 186.300 152.700 186.700 152.800 ;
        RECT 186.300 152.400 187.700 152.700 ;
        RECT 187.400 152.100 187.700 152.400 ;
        RECT 189.400 152.100 189.800 152.500 ;
        RECT 184.600 151.800 185.600 152.100 ;
        RECT 185.200 151.100 185.600 151.800 ;
        RECT 187.400 151.100 187.800 152.100 ;
        RECT 189.400 151.800 190.100 152.100 ;
        RECT 189.500 151.100 190.100 151.800 ;
        RECT 191.800 151.100 192.200 153.300 ;
        RECT 192.600 153.400 193.700 153.700 ;
        RECT 192.600 151.100 193.000 153.400 ;
        RECT 0.600 147.700 1.000 149.900 ;
        RECT 2.700 149.200 3.300 149.900 ;
        RECT 2.700 148.900 3.400 149.200 ;
        RECT 5.000 148.900 5.400 149.900 ;
        RECT 7.200 149.200 7.600 149.900 ;
        RECT 7.200 148.900 8.200 149.200 ;
        RECT 3.000 148.500 3.400 148.900 ;
        RECT 5.100 148.600 5.400 148.900 ;
        RECT 5.100 148.300 6.500 148.600 ;
        RECT 6.100 148.200 6.500 148.300 ;
        RECT 7.000 148.200 7.400 148.600 ;
        RECT 7.800 148.500 8.200 148.900 ;
        RECT 2.100 147.700 2.500 147.800 ;
        RECT 0.600 147.400 2.500 147.700 ;
        RECT 0.600 145.700 1.000 147.400 ;
        RECT 4.100 147.100 4.500 147.200 ;
        RECT 7.000 147.100 7.300 148.200 ;
        RECT 9.400 147.500 9.800 149.900 ;
        RECT 11.000 148.900 11.400 149.900 ;
        RECT 10.200 147.800 10.600 148.600 ;
        RECT 8.600 147.100 9.400 147.200 ;
        RECT 10.200 147.100 10.500 147.800 ;
        RECT 11.100 147.200 11.400 148.900 ;
        RECT 3.900 146.800 10.500 147.100 ;
        RECT 11.000 146.800 11.400 147.200 ;
        RECT 12.600 148.500 13.000 149.500 ;
        RECT 12.600 147.400 12.900 148.500 ;
        RECT 14.700 148.000 15.100 149.500 ;
        RECT 14.700 147.700 15.500 148.000 ;
        RECT 15.100 147.500 15.500 147.700 ;
        RECT 12.600 147.100 14.700 147.400 ;
        RECT 3.000 146.400 3.400 146.500 ;
        RECT 1.500 146.100 3.400 146.400 ;
        RECT 1.500 146.000 1.900 146.100 ;
        RECT 2.300 145.700 2.700 145.800 ;
        RECT 0.600 145.400 2.700 145.700 ;
        RECT 0.600 141.100 1.000 145.400 ;
        RECT 3.900 145.200 4.200 146.800 ;
        RECT 7.500 146.700 7.900 146.800 ;
        RECT 8.300 146.200 8.700 146.300 ;
        RECT 11.100 146.200 11.400 146.800 ;
        RECT 14.200 146.900 14.700 147.100 ;
        RECT 15.200 147.200 15.500 147.500 ;
        RECT 17.400 147.700 17.800 149.900 ;
        RECT 19.500 149.200 20.100 149.900 ;
        RECT 19.500 148.900 20.200 149.200 ;
        RECT 21.800 148.900 22.200 149.900 ;
        RECT 24.000 149.200 24.400 149.900 ;
        RECT 24.000 148.900 25.000 149.200 ;
        RECT 19.800 148.500 20.200 148.900 ;
        RECT 21.900 148.600 22.200 148.900 ;
        RECT 21.900 148.300 23.300 148.600 ;
        RECT 22.900 148.200 23.300 148.300 ;
        RECT 23.800 148.200 24.200 148.600 ;
        RECT 24.600 148.500 25.000 148.900 ;
        RECT 18.900 147.700 19.300 147.800 ;
        RECT 17.400 147.400 19.300 147.700 ;
        RECT 6.200 145.900 8.700 146.200 ;
        RECT 6.200 145.800 6.600 145.900 ;
        RECT 11.000 145.800 11.400 146.200 ;
        RECT 7.000 145.500 9.800 145.600 ;
        RECT 6.900 145.400 9.800 145.500 ;
        RECT 3.000 144.900 4.200 145.200 ;
        RECT 4.900 145.300 9.800 145.400 ;
        RECT 4.900 145.100 7.300 145.300 ;
        RECT 3.000 144.400 3.300 144.900 ;
        RECT 2.600 144.000 3.300 144.400 ;
        RECT 4.100 144.500 4.500 144.600 ;
        RECT 4.900 144.500 5.200 145.100 ;
        RECT 4.100 144.200 5.200 144.500 ;
        RECT 5.500 144.500 8.200 144.800 ;
        RECT 5.500 144.400 5.900 144.500 ;
        RECT 7.800 144.400 8.200 144.500 ;
        RECT 4.700 143.700 5.100 143.800 ;
        RECT 6.100 143.700 6.500 143.800 ;
        RECT 3.000 143.100 3.400 143.500 ;
        RECT 4.700 143.400 6.500 143.700 ;
        RECT 5.100 143.100 5.400 143.400 ;
        RECT 7.800 143.100 8.200 143.500 ;
        RECT 2.700 141.100 3.300 143.100 ;
        RECT 5.000 141.100 5.400 143.100 ;
        RECT 7.200 142.800 8.200 143.100 ;
        RECT 7.200 141.100 7.600 142.800 ;
        RECT 9.400 141.100 9.800 145.300 ;
        RECT 11.100 145.100 11.400 145.800 ;
        RECT 11.800 145.400 12.200 146.200 ;
        RECT 12.600 145.800 13.000 146.600 ;
        RECT 13.400 145.800 13.800 146.600 ;
        RECT 14.200 146.500 14.900 146.900 ;
        RECT 15.200 146.800 16.200 147.200 ;
        RECT 14.200 145.500 14.500 146.500 ;
        RECT 15.200 146.200 15.500 146.800 ;
        RECT 15.000 145.800 15.500 146.200 ;
        RECT 12.600 145.200 14.500 145.500 ;
        RECT 11.000 144.700 11.900 145.100 ;
        RECT 11.500 141.100 11.900 144.700 ;
        RECT 12.600 143.500 12.900 145.200 ;
        RECT 15.200 144.900 15.500 145.800 ;
        RECT 15.800 146.100 16.200 146.200 ;
        RECT 16.600 146.100 17.000 146.200 ;
        RECT 15.800 145.800 17.000 146.100 ;
        RECT 15.800 145.400 16.200 145.800 ;
        RECT 17.400 145.700 17.800 147.400 ;
        RECT 20.900 147.100 21.300 147.200 ;
        RECT 23.800 147.100 24.100 148.200 ;
        RECT 26.200 147.500 26.600 149.900 ;
        RECT 27.000 147.700 27.400 149.900 ;
        RECT 29.100 149.200 29.700 149.900 ;
        RECT 29.100 148.900 29.800 149.200 ;
        RECT 31.400 148.900 31.800 149.900 ;
        RECT 33.600 149.200 34.000 149.900 ;
        RECT 33.600 148.900 34.600 149.200 ;
        RECT 29.400 148.500 29.800 148.900 ;
        RECT 31.500 148.600 31.800 148.900 ;
        RECT 31.500 148.300 32.900 148.600 ;
        RECT 32.500 148.200 32.900 148.300 ;
        RECT 33.400 148.200 33.800 148.600 ;
        RECT 34.200 148.500 34.600 148.900 ;
        RECT 28.500 147.700 28.900 147.800 ;
        RECT 27.000 147.400 28.900 147.700 ;
        RECT 25.400 147.100 26.200 147.200 ;
        RECT 20.700 146.800 26.200 147.100 ;
        RECT 19.800 146.400 20.200 146.500 ;
        RECT 18.300 146.100 20.200 146.400 ;
        RECT 20.700 146.200 21.000 146.800 ;
        RECT 24.300 146.700 24.700 146.800 ;
        RECT 23.800 146.200 24.200 146.300 ;
        RECT 25.100 146.200 25.500 146.300 ;
        RECT 18.300 146.000 18.700 146.100 ;
        RECT 20.600 145.800 21.000 146.200 ;
        RECT 23.000 145.900 25.500 146.200 ;
        RECT 23.000 145.800 23.400 145.900 ;
        RECT 19.100 145.700 19.500 145.800 ;
        RECT 17.400 145.400 19.500 145.700 ;
        RECT 14.700 144.600 15.500 144.900 ;
        RECT 12.600 141.500 13.000 143.500 ;
        RECT 14.700 141.100 15.100 144.600 ;
        RECT 17.400 141.100 17.800 145.400 ;
        RECT 20.700 145.200 21.000 145.800 ;
        RECT 27.000 145.700 27.400 147.400 ;
        RECT 30.500 147.100 30.900 147.200 ;
        RECT 32.600 147.100 33.000 147.200 ;
        RECT 33.400 147.100 33.700 148.200 ;
        RECT 35.800 147.500 36.200 149.900 ;
        RECT 36.600 147.900 37.000 149.900 ;
        RECT 37.400 148.000 37.800 149.900 ;
        RECT 39.000 148.000 39.400 149.900 ;
        RECT 39.900 148.200 40.300 148.600 ;
        RECT 37.400 147.900 39.400 148.000 ;
        RECT 36.700 147.200 37.000 147.900 ;
        RECT 37.500 147.700 39.300 147.900 ;
        RECT 39.800 147.800 40.200 148.200 ;
        RECT 40.600 147.900 41.000 149.900 ;
        RECT 38.600 147.200 39.000 147.400 ;
        RECT 35.000 147.100 35.800 147.200 ;
        RECT 30.300 146.800 35.800 147.100 ;
        RECT 36.600 146.800 37.900 147.200 ;
        RECT 38.600 146.900 39.400 147.200 ;
        RECT 39.000 146.800 39.400 146.900 ;
        RECT 29.400 146.400 29.800 146.500 ;
        RECT 27.900 146.100 29.800 146.400 ;
        RECT 27.900 146.000 28.300 146.100 ;
        RECT 28.700 145.700 29.100 145.800 ;
        RECT 23.800 145.500 26.600 145.600 ;
        RECT 23.700 145.400 26.600 145.500 ;
        RECT 19.800 144.900 21.000 145.200 ;
        RECT 21.700 145.300 26.600 145.400 ;
        RECT 21.700 145.100 24.100 145.300 ;
        RECT 19.800 144.400 20.100 144.900 ;
        RECT 19.400 144.000 20.100 144.400 ;
        RECT 20.900 144.500 21.300 144.600 ;
        RECT 21.700 144.500 22.000 145.100 ;
        RECT 20.900 144.200 22.000 144.500 ;
        RECT 22.300 144.500 25.000 144.800 ;
        RECT 22.300 144.400 22.700 144.500 ;
        RECT 24.600 144.400 25.000 144.500 ;
        RECT 21.500 143.700 21.900 143.800 ;
        RECT 22.900 143.700 23.300 143.800 ;
        RECT 19.800 143.100 20.200 143.500 ;
        RECT 21.500 143.400 23.300 143.700 ;
        RECT 21.900 143.100 22.200 143.400 ;
        RECT 24.600 143.100 25.000 143.500 ;
        RECT 19.500 141.100 20.100 143.100 ;
        RECT 21.800 141.100 22.200 143.100 ;
        RECT 24.000 142.800 25.000 143.100 ;
        RECT 24.000 141.100 24.400 142.800 ;
        RECT 26.200 141.100 26.600 145.300 ;
        RECT 27.000 145.400 29.100 145.700 ;
        RECT 27.000 141.100 27.400 145.400 ;
        RECT 30.300 145.200 30.600 146.800 ;
        RECT 33.900 146.700 34.300 146.800 ;
        RECT 33.400 146.200 33.800 146.300 ;
        RECT 34.700 146.200 35.100 146.300 ;
        RECT 32.600 145.900 35.100 146.200 ;
        RECT 32.600 145.800 33.000 145.900 ;
        RECT 33.400 145.500 36.200 145.600 ;
        RECT 33.300 145.400 36.200 145.500 ;
        RECT 29.400 144.900 30.600 145.200 ;
        RECT 31.300 145.300 36.200 145.400 ;
        RECT 31.300 145.100 33.700 145.300 ;
        RECT 29.400 144.400 29.700 144.900 ;
        RECT 29.000 144.200 29.700 144.400 ;
        RECT 30.500 144.500 30.900 144.600 ;
        RECT 31.300 144.500 31.600 145.100 ;
        RECT 30.500 144.200 31.600 144.500 ;
        RECT 31.900 144.500 34.600 144.800 ;
        RECT 31.900 144.400 32.300 144.500 ;
        RECT 34.200 144.400 34.600 144.500 ;
        RECT 28.600 144.000 29.700 144.200 ;
        RECT 28.600 143.800 29.300 144.000 ;
        RECT 31.100 143.700 31.500 143.800 ;
        RECT 32.500 143.700 32.900 143.800 ;
        RECT 29.400 143.100 29.800 143.500 ;
        RECT 31.100 143.400 32.900 143.700 ;
        RECT 31.500 143.100 31.800 143.400 ;
        RECT 34.200 143.100 34.600 143.500 ;
        RECT 29.100 141.100 29.700 143.100 ;
        RECT 31.400 141.100 31.800 143.100 ;
        RECT 33.600 142.800 34.600 143.100 ;
        RECT 33.600 141.100 34.000 142.800 ;
        RECT 35.800 141.100 36.200 145.300 ;
        RECT 36.600 145.100 37.000 145.200 ;
        RECT 37.600 145.100 37.900 146.800 ;
        RECT 38.200 145.800 38.600 146.600 ;
        RECT 39.800 146.100 40.200 146.200 ;
        RECT 40.700 146.100 41.000 147.900 ;
        RECT 41.400 146.400 41.800 147.200 ;
        RECT 43.000 146.800 43.400 147.600 ;
        RECT 43.800 147.100 44.200 149.900 ;
        RECT 46.200 147.900 46.600 149.900 ;
        RECT 48.400 148.100 49.200 149.900 ;
        RECT 46.200 147.600 47.400 147.900 ;
        RECT 47.000 147.500 47.400 147.600 ;
        RECT 47.700 147.400 48.100 147.800 ;
        RECT 47.700 147.200 48.000 147.400 ;
        RECT 46.200 147.100 47.000 147.200 ;
        RECT 43.800 146.800 47.000 147.100 ;
        RECT 47.600 146.800 48.000 147.200 ;
        RECT 42.200 146.100 42.600 146.200 ;
        RECT 39.800 145.800 41.000 146.100 ;
        RECT 41.800 145.800 42.600 146.100 ;
        RECT 39.900 145.100 40.200 145.800 ;
        RECT 41.800 145.600 42.200 145.800 ;
        RECT 36.600 144.800 37.300 145.100 ;
        RECT 37.600 144.800 38.100 145.100 ;
        RECT 37.000 144.200 37.300 144.800 ;
        RECT 37.000 143.800 37.400 144.200 ;
        RECT 37.700 141.100 38.100 144.800 ;
        RECT 39.800 141.100 40.200 145.100 ;
        RECT 40.600 144.800 42.600 145.100 ;
        RECT 40.600 141.100 41.000 144.800 ;
        RECT 42.200 141.100 42.600 144.800 ;
        RECT 43.800 141.100 44.200 146.800 ;
        RECT 48.400 146.400 48.700 148.100 ;
        RECT 51.000 147.900 51.400 149.900 ;
        RECT 49.000 147.700 49.800 147.800 ;
        RECT 49.000 147.400 50.000 147.700 ;
        RECT 50.300 147.600 51.400 147.900 ;
        RECT 53.400 147.800 53.800 149.900 ;
        RECT 54.100 148.200 54.500 148.600 ;
        RECT 54.200 148.100 54.600 148.200 ;
        RECT 55.000 148.100 55.400 149.900 ;
        RECT 54.200 147.800 55.400 148.100 ;
        RECT 55.800 148.000 56.200 149.900 ;
        RECT 57.400 148.000 57.800 149.900 ;
        RECT 55.800 147.900 57.800 148.000 ;
        RECT 50.300 147.500 50.700 147.600 ;
        RECT 49.700 147.200 50.000 147.400 ;
        RECT 49.000 146.700 49.400 147.100 ;
        RECT 49.700 146.900 51.400 147.200 ;
        RECT 50.600 146.800 51.400 146.900 ;
        RECT 48.200 146.200 48.700 146.400 ;
        RECT 45.400 146.100 45.800 146.200 ;
        RECT 47.800 146.100 48.700 146.200 ;
        RECT 49.100 146.400 49.400 146.700 ;
        RECT 52.600 146.400 53.000 147.200 ;
        RECT 49.100 146.100 50.400 146.400 ;
        RECT 45.400 145.800 48.500 146.100 ;
        RECT 50.000 146.000 50.400 146.100 ;
        RECT 51.800 146.100 52.200 146.200 ;
        RECT 53.400 146.100 53.700 147.800 ;
        RECT 55.100 147.200 55.400 147.800 ;
        RECT 55.900 147.700 57.700 147.900 ;
        RECT 57.000 147.200 57.400 147.400 ;
        RECT 55.000 146.800 56.300 147.200 ;
        RECT 57.000 146.900 57.800 147.200 ;
        RECT 57.400 146.800 57.800 146.900 ;
        RECT 58.200 146.800 58.600 147.600 ;
        RECT 54.200 146.100 54.600 146.200 ;
        RECT 51.800 145.800 52.600 146.100 ;
        RECT 53.400 145.800 54.600 146.100 ;
        RECT 48.200 145.100 48.500 145.800 ;
        RECT 48.900 145.700 49.300 145.800 ;
        RECT 48.900 145.400 50.600 145.700 ;
        RECT 52.200 145.600 52.600 145.800 ;
        RECT 50.300 145.100 50.600 145.400 ;
        RECT 54.200 145.100 54.500 145.800 ;
        RECT 55.000 145.100 55.400 145.200 ;
        RECT 56.000 145.100 56.300 146.800 ;
        RECT 56.600 145.800 57.000 146.600 ;
        RECT 46.200 144.800 47.400 145.100 ;
        RECT 48.200 144.800 49.200 145.100 ;
        RECT 46.200 141.100 46.600 144.800 ;
        RECT 47.000 144.700 47.400 144.800 ;
        RECT 48.400 141.100 49.200 144.800 ;
        RECT 50.300 144.800 51.400 145.100 ;
        RECT 50.300 144.700 50.700 144.800 ;
        RECT 51.000 141.100 51.400 144.800 ;
        RECT 51.800 144.800 53.800 145.100 ;
        RECT 51.800 141.100 52.200 144.800 ;
        RECT 53.400 141.100 53.800 144.800 ;
        RECT 54.200 141.100 54.600 145.100 ;
        RECT 55.000 144.800 55.700 145.100 ;
        RECT 56.000 144.800 56.500 145.100 ;
        RECT 55.400 144.200 55.700 144.800 ;
        RECT 55.400 143.800 55.800 144.200 ;
        RECT 56.100 141.100 56.500 144.800 ;
        RECT 59.000 141.100 59.400 149.900 ;
        RECT 61.400 147.900 61.800 149.900 ;
        RECT 62.100 148.200 62.500 148.600 ;
        RECT 63.000 148.500 63.400 149.500 ;
        RECT 65.100 149.200 65.500 149.500 ;
        RECT 64.600 148.800 65.500 149.200 ;
        RECT 60.600 146.400 61.000 147.200 ;
        RECT 59.800 146.100 60.200 146.200 ;
        RECT 61.400 146.100 61.700 147.900 ;
        RECT 62.200 147.800 62.600 148.200 ;
        RECT 63.000 147.400 63.300 148.500 ;
        RECT 65.100 148.000 65.500 148.800 ;
        RECT 68.600 148.200 69.000 149.900 ;
        RECT 65.100 147.700 65.900 148.000 ;
        RECT 65.500 147.500 65.900 147.700 ;
        RECT 63.000 147.100 65.100 147.400 ;
        RECT 64.600 146.900 65.100 147.100 ;
        RECT 65.600 147.200 65.900 147.500 ;
        RECT 68.500 147.900 69.000 148.200 ;
        RECT 68.500 147.200 68.800 147.900 ;
        RECT 70.200 147.600 70.600 149.900 ;
        RECT 71.000 147.800 71.400 149.900 ;
        RECT 71.800 148.000 72.200 149.900 ;
        RECT 73.400 148.000 73.800 149.900 ;
        RECT 71.800 147.900 73.800 148.000 ;
        RECT 69.300 147.300 70.600 147.600 ;
        RECT 62.200 146.100 62.600 146.200 ;
        RECT 59.800 145.800 60.600 146.100 ;
        RECT 61.400 145.800 62.600 146.100 ;
        RECT 63.000 145.800 63.400 146.600 ;
        RECT 63.800 145.800 64.200 146.600 ;
        RECT 64.600 146.500 65.300 146.900 ;
        RECT 65.600 146.800 66.600 147.200 ;
        RECT 68.500 146.800 69.000 147.200 ;
        RECT 60.200 145.600 60.600 145.800 ;
        RECT 62.200 145.100 62.500 145.800 ;
        RECT 64.600 145.500 64.900 146.500 ;
        RECT 63.000 145.200 64.900 145.500 ;
        RECT 59.800 144.800 61.800 145.100 ;
        RECT 59.800 141.100 60.200 144.800 ;
        RECT 61.400 141.100 61.800 144.800 ;
        RECT 62.200 141.100 62.600 145.100 ;
        RECT 63.000 143.500 63.300 145.200 ;
        RECT 65.600 144.900 65.900 146.800 ;
        RECT 66.200 145.400 66.600 146.200 ;
        RECT 65.100 144.600 65.900 144.900 ;
        RECT 68.500 145.100 68.800 146.800 ;
        RECT 69.300 146.500 69.600 147.300 ;
        RECT 71.100 147.200 71.400 147.800 ;
        RECT 71.900 147.700 73.700 147.900 ;
        RECT 74.200 147.700 74.600 149.900 ;
        RECT 76.300 149.200 76.900 149.900 ;
        RECT 76.300 148.900 77.000 149.200 ;
        RECT 78.600 148.900 79.000 149.900 ;
        RECT 80.800 149.200 81.200 149.900 ;
        RECT 80.800 148.900 81.800 149.200 ;
        RECT 76.600 148.500 77.000 148.900 ;
        RECT 78.700 148.600 79.000 148.900 ;
        RECT 78.700 148.300 80.100 148.600 ;
        RECT 79.700 148.200 80.100 148.300 ;
        RECT 80.600 148.200 81.000 148.600 ;
        RECT 81.400 148.500 81.800 148.900 ;
        RECT 75.700 147.700 76.100 147.800 ;
        RECT 74.200 147.400 76.100 147.700 ;
        RECT 73.000 147.200 73.400 147.400 ;
        RECT 71.000 146.800 72.300 147.200 ;
        RECT 73.000 146.900 73.800 147.200 ;
        RECT 73.400 146.800 73.800 146.900 ;
        RECT 69.100 146.100 69.600 146.500 ;
        RECT 69.300 145.100 69.600 146.100 ;
        RECT 70.100 146.200 70.500 146.600 ;
        RECT 70.100 145.800 70.600 146.200 ;
        RECT 71.000 145.100 71.400 145.200 ;
        RECT 72.000 145.100 72.300 146.800 ;
        RECT 72.600 146.100 73.000 146.600 ;
        RECT 74.200 146.100 74.600 147.400 ;
        RECT 77.400 147.100 78.100 147.200 ;
        RECT 80.600 147.100 80.900 148.200 ;
        RECT 83.000 147.500 83.400 149.900 ;
        RECT 84.600 148.900 85.000 149.900 ;
        RECT 83.800 147.800 84.200 148.600 ;
        RECT 84.700 147.200 85.000 148.900 ;
        RECT 87.800 147.900 88.200 149.900 ;
        RECT 88.500 148.200 88.900 148.600 ;
        RECT 88.600 148.100 89.000 148.200 ;
        RECT 89.400 148.100 89.800 149.900 ;
        RECT 82.200 147.100 83.000 147.200 ;
        RECT 77.400 146.800 83.000 147.100 ;
        RECT 83.800 146.800 84.200 147.200 ;
        RECT 84.600 146.800 85.000 147.200 ;
        RECT 76.600 146.400 77.000 146.500 ;
        RECT 72.600 145.800 74.600 146.100 ;
        RECT 75.100 146.100 77.000 146.400 ;
        RECT 75.100 146.000 75.500 146.100 ;
        RECT 74.200 145.700 74.600 145.800 ;
        RECT 75.900 145.700 76.300 145.800 ;
        RECT 74.200 145.400 76.300 145.700 ;
        RECT 68.500 144.600 69.000 145.100 ;
        RECT 69.300 144.800 70.600 145.100 ;
        RECT 71.000 144.800 71.700 145.100 ;
        RECT 72.000 144.800 72.500 145.100 ;
        RECT 63.000 141.500 63.400 143.500 ;
        RECT 65.100 141.100 65.500 144.600 ;
        RECT 68.600 141.100 69.000 144.600 ;
        RECT 70.200 141.100 70.600 144.800 ;
        RECT 71.400 144.200 71.700 144.800 ;
        RECT 71.400 143.800 71.800 144.200 ;
        RECT 72.100 141.100 72.500 144.800 ;
        RECT 74.200 141.100 74.600 145.400 ;
        RECT 77.500 145.200 77.800 146.800 ;
        RECT 81.100 146.700 81.500 146.800 ;
        RECT 80.600 146.200 81.000 146.300 ;
        RECT 81.900 146.200 82.300 146.300 ;
        RECT 79.800 145.900 82.300 146.200 ;
        RECT 83.800 146.100 84.100 146.800 ;
        RECT 84.700 146.100 85.000 146.800 ;
        RECT 87.000 146.400 87.400 147.200 ;
        RECT 79.800 145.800 80.200 145.900 ;
        RECT 83.800 145.800 85.000 146.100 ;
        RECT 80.600 145.500 83.400 145.600 ;
        RECT 80.500 145.400 83.400 145.500 ;
        RECT 76.600 144.900 77.800 145.200 ;
        RECT 78.500 145.300 83.400 145.400 ;
        RECT 78.500 145.100 80.900 145.300 ;
        RECT 76.600 144.400 76.900 144.900 ;
        RECT 76.200 144.000 76.900 144.400 ;
        RECT 77.700 144.500 78.100 144.600 ;
        RECT 78.500 144.500 78.800 145.100 ;
        RECT 77.700 144.200 78.800 144.500 ;
        RECT 79.100 144.500 81.800 144.800 ;
        RECT 79.100 144.400 79.500 144.500 ;
        RECT 81.400 144.400 81.800 144.500 ;
        RECT 78.300 143.700 78.700 143.800 ;
        RECT 79.700 143.700 80.100 143.800 ;
        RECT 76.600 143.100 77.000 143.500 ;
        RECT 78.300 143.400 80.100 143.700 ;
        RECT 78.700 143.100 79.000 143.400 ;
        RECT 81.400 143.100 81.800 143.500 ;
        RECT 76.300 141.100 76.900 143.100 ;
        RECT 78.600 141.100 79.000 143.100 ;
        RECT 80.800 142.800 81.800 143.100 ;
        RECT 80.800 141.100 81.200 142.800 ;
        RECT 83.000 141.100 83.400 145.300 ;
        RECT 84.700 145.100 85.000 145.800 ;
        RECT 85.400 145.400 85.800 146.200 ;
        RECT 86.200 146.100 86.600 146.200 ;
        RECT 87.800 146.100 88.100 147.900 ;
        RECT 88.600 147.800 89.800 148.100 ;
        RECT 90.200 148.000 90.600 149.900 ;
        RECT 91.800 148.000 92.200 149.900 ;
        RECT 94.500 149.200 94.900 149.500 ;
        RECT 94.500 148.800 95.400 149.200 ;
        RECT 94.500 148.000 94.900 148.800 ;
        RECT 96.600 148.500 97.000 149.500 ;
        RECT 90.200 147.900 92.200 148.000 ;
        RECT 89.500 147.200 89.800 147.800 ;
        RECT 90.300 147.700 92.100 147.900 ;
        RECT 94.100 147.700 94.900 148.000 ;
        RECT 94.100 147.500 94.500 147.700 ;
        RECT 91.400 147.200 91.800 147.400 ;
        RECT 94.100 147.200 94.400 147.500 ;
        RECT 96.700 147.400 97.000 148.500 ;
        RECT 89.400 146.800 90.700 147.200 ;
        RECT 91.400 146.900 92.200 147.200 ;
        RECT 91.800 146.800 92.200 146.900 ;
        RECT 93.400 146.800 94.400 147.200 ;
        RECT 94.900 147.100 97.000 147.400 ;
        RECT 99.000 148.500 99.400 149.500 ;
        RECT 101.100 149.200 101.500 149.500 ;
        RECT 101.100 148.800 101.800 149.200 ;
        RECT 99.000 147.400 99.300 148.500 ;
        RECT 101.100 148.000 101.500 148.800 ;
        RECT 101.100 147.700 101.900 148.000 ;
        RECT 101.500 147.500 101.900 147.700 ;
        RECT 99.000 147.100 101.100 147.400 ;
        RECT 94.900 146.900 95.400 147.100 ;
        RECT 88.600 146.100 89.000 146.200 ;
        RECT 86.200 145.800 87.000 146.100 ;
        RECT 87.800 145.800 89.000 146.100 ;
        RECT 86.600 145.600 87.000 145.800 ;
        RECT 88.600 145.100 88.900 145.800 ;
        RECT 89.400 145.100 89.800 145.200 ;
        RECT 90.400 145.100 90.700 146.800 ;
        RECT 91.000 145.800 91.400 146.600 ;
        RECT 93.400 145.400 93.800 146.200 ;
        RECT 84.600 144.700 85.500 145.100 ;
        RECT 85.100 141.100 85.500 144.700 ;
        RECT 86.200 144.800 88.200 145.100 ;
        RECT 86.200 141.100 86.600 144.800 ;
        RECT 87.800 141.100 88.200 144.800 ;
        RECT 88.600 141.100 89.000 145.100 ;
        RECT 89.400 144.800 90.100 145.100 ;
        RECT 90.400 144.800 90.900 145.100 ;
        RECT 89.800 144.200 90.100 144.800 ;
        RECT 89.800 143.800 90.200 144.200 ;
        RECT 90.500 141.100 90.900 144.800 ;
        RECT 94.100 144.900 94.400 146.800 ;
        RECT 94.700 146.500 95.400 146.900 ;
        RECT 100.600 146.900 101.100 147.100 ;
        RECT 101.600 147.200 101.900 147.500 ;
        RECT 103.800 147.700 104.200 149.900 ;
        RECT 105.900 149.200 106.500 149.900 ;
        RECT 105.900 148.900 106.600 149.200 ;
        RECT 108.200 148.900 108.600 149.900 ;
        RECT 110.400 149.200 110.800 149.900 ;
        RECT 110.400 148.900 111.400 149.200 ;
        RECT 106.200 148.500 106.600 148.900 ;
        RECT 108.300 148.600 108.600 148.900 ;
        RECT 108.300 148.300 109.700 148.600 ;
        RECT 109.300 148.200 109.700 148.300 ;
        RECT 110.200 148.200 110.600 148.600 ;
        RECT 111.000 148.500 111.400 148.900 ;
        RECT 105.300 147.700 105.700 147.800 ;
        RECT 103.800 147.400 105.700 147.700 ;
        RECT 95.100 145.500 95.400 146.500 ;
        RECT 95.800 145.800 96.200 146.600 ;
        RECT 96.600 146.100 97.000 146.600 ;
        RECT 99.000 146.100 99.400 146.600 ;
        RECT 96.600 145.800 99.400 146.100 ;
        RECT 99.800 145.800 100.200 146.600 ;
        RECT 100.600 146.500 101.300 146.900 ;
        RECT 101.600 146.800 102.600 147.200 ;
        RECT 100.600 145.500 100.900 146.500 ;
        RECT 95.100 145.200 97.000 145.500 ;
        RECT 94.100 144.600 94.900 144.900 ;
        RECT 94.500 141.100 94.900 144.600 ;
        RECT 96.700 143.500 97.000 145.200 ;
        RECT 96.600 141.500 97.000 143.500 ;
        RECT 99.000 145.200 100.900 145.500 ;
        RECT 99.000 143.500 99.300 145.200 ;
        RECT 101.600 144.900 101.900 146.800 ;
        RECT 102.200 146.100 102.600 146.200 ;
        RECT 103.800 146.100 104.200 147.400 ;
        RECT 107.300 147.100 107.700 147.200 ;
        RECT 110.200 147.100 110.500 148.200 ;
        RECT 112.600 147.500 113.000 149.900 ;
        RECT 113.400 147.700 113.800 149.900 ;
        RECT 115.500 149.200 116.100 149.900 ;
        RECT 115.500 148.900 116.200 149.200 ;
        RECT 117.800 148.900 118.200 149.900 ;
        RECT 120.000 149.200 120.400 149.900 ;
        RECT 120.000 148.900 121.000 149.200 ;
        RECT 115.800 148.500 116.200 148.900 ;
        RECT 117.900 148.600 118.200 148.900 ;
        RECT 117.900 148.300 119.300 148.600 ;
        RECT 118.900 148.200 119.300 148.300 ;
        RECT 119.800 148.200 120.200 148.600 ;
        RECT 120.600 148.500 121.000 148.900 ;
        RECT 114.900 147.700 115.300 147.800 ;
        RECT 113.400 147.400 115.300 147.700 ;
        RECT 111.800 147.100 112.600 147.200 ;
        RECT 107.100 146.800 112.600 147.100 ;
        RECT 106.200 146.400 106.600 146.500 ;
        RECT 102.200 145.800 104.200 146.100 ;
        RECT 104.700 146.100 106.600 146.400 ;
        RECT 107.100 146.200 107.400 146.800 ;
        RECT 110.700 146.700 111.100 146.800 ;
        RECT 110.200 146.200 110.600 146.300 ;
        RECT 111.500 146.200 111.900 146.300 ;
        RECT 104.700 146.000 105.100 146.100 ;
        RECT 107.000 145.800 107.400 146.200 ;
        RECT 109.400 145.900 111.900 146.200 ;
        RECT 109.400 145.800 109.800 145.900 ;
        RECT 102.200 145.400 102.600 145.800 ;
        RECT 103.800 145.700 104.200 145.800 ;
        RECT 105.500 145.700 105.900 145.800 ;
        RECT 103.800 145.400 105.900 145.700 ;
        RECT 101.100 144.600 101.900 144.900 ;
        RECT 99.000 141.500 99.400 143.500 ;
        RECT 101.100 141.100 101.500 144.600 ;
        RECT 103.800 141.100 104.200 145.400 ;
        RECT 107.100 145.200 107.400 145.800 ;
        RECT 113.400 145.700 113.800 147.400 ;
        RECT 116.900 147.100 117.300 147.200 ;
        RECT 119.800 147.100 120.100 148.200 ;
        RECT 122.200 147.500 122.600 149.900 ;
        RECT 123.800 148.900 124.200 149.900 ;
        RECT 123.000 148.100 123.400 148.200 ;
        RECT 123.800 148.100 124.100 148.900 ;
        RECT 123.000 147.800 124.100 148.100 ;
        RECT 124.600 147.800 125.000 148.600 ;
        RECT 123.800 147.200 124.100 147.800 ;
        RECT 126.200 147.600 126.600 149.900 ;
        RECT 127.800 147.600 128.200 149.900 ;
        RECT 129.400 147.600 129.800 149.900 ;
        RECT 131.000 147.600 131.400 149.900 ;
        RECT 125.400 147.200 126.600 147.600 ;
        RECT 127.100 147.200 128.200 147.600 ;
        RECT 128.700 147.200 129.800 147.600 ;
        RECT 130.500 147.200 131.400 147.600 ;
        RECT 132.600 147.700 133.000 149.900 ;
        RECT 134.700 149.200 135.300 149.900 ;
        RECT 134.700 148.900 135.400 149.200 ;
        RECT 137.000 148.900 137.400 149.900 ;
        RECT 139.200 149.200 139.600 149.900 ;
        RECT 139.200 148.900 140.200 149.200 ;
        RECT 135.000 148.500 135.400 148.900 ;
        RECT 137.100 148.600 137.400 148.900 ;
        RECT 137.100 148.300 138.500 148.600 ;
        RECT 138.100 148.200 138.500 148.300 ;
        RECT 139.000 148.200 139.400 148.600 ;
        RECT 139.800 148.500 140.200 148.900 ;
        RECT 134.100 147.700 134.500 147.800 ;
        RECT 132.600 147.400 134.500 147.700 ;
        RECT 121.400 147.100 122.200 147.200 ;
        RECT 116.700 146.800 122.200 147.100 ;
        RECT 123.800 146.800 124.200 147.200 ;
        RECT 115.800 146.400 116.200 146.500 ;
        RECT 114.300 146.100 116.200 146.400 ;
        RECT 114.300 146.000 114.700 146.100 ;
        RECT 115.100 145.700 115.500 145.800 ;
        RECT 110.200 145.500 113.000 145.600 ;
        RECT 110.100 145.400 113.000 145.500 ;
        RECT 106.200 144.900 107.400 145.200 ;
        RECT 108.100 145.300 113.000 145.400 ;
        RECT 108.100 145.100 110.500 145.300 ;
        RECT 106.200 144.400 106.500 144.900 ;
        RECT 105.800 144.000 106.500 144.400 ;
        RECT 107.300 144.500 107.700 144.600 ;
        RECT 108.100 144.500 108.400 145.100 ;
        RECT 107.300 144.200 108.400 144.500 ;
        RECT 108.700 144.500 111.400 144.800 ;
        RECT 108.700 144.400 109.100 144.500 ;
        RECT 111.000 144.400 111.400 144.500 ;
        RECT 107.900 143.700 108.300 143.800 ;
        RECT 109.300 143.700 109.700 143.800 ;
        RECT 106.200 143.100 106.600 143.500 ;
        RECT 107.900 143.400 109.700 143.700 ;
        RECT 108.300 143.100 108.600 143.400 ;
        RECT 111.000 143.100 111.400 143.500 ;
        RECT 105.900 141.100 106.500 143.100 ;
        RECT 108.200 141.100 108.600 143.100 ;
        RECT 110.400 142.800 111.400 143.100 ;
        RECT 110.400 141.100 110.800 142.800 ;
        RECT 112.600 141.100 113.000 145.300 ;
        RECT 113.400 145.400 115.500 145.700 ;
        RECT 113.400 141.100 113.800 145.400 ;
        RECT 116.700 145.200 117.000 146.800 ;
        RECT 120.300 146.700 120.700 146.800 ;
        RECT 119.800 146.200 120.200 146.300 ;
        RECT 121.100 146.200 121.500 146.300 ;
        RECT 119.000 145.900 121.500 146.200 ;
        RECT 119.000 145.800 119.400 145.900 ;
        RECT 119.800 145.500 122.600 145.600 ;
        RECT 119.700 145.400 122.600 145.500 ;
        RECT 123.000 145.400 123.400 146.200 ;
        RECT 115.800 144.900 117.000 145.200 ;
        RECT 117.700 145.300 122.600 145.400 ;
        RECT 117.700 145.100 120.100 145.300 ;
        RECT 115.800 144.400 116.100 144.900 ;
        RECT 115.400 144.000 116.100 144.400 ;
        RECT 116.900 144.500 117.300 144.600 ;
        RECT 117.700 144.500 118.000 145.100 ;
        RECT 116.900 144.200 118.000 144.500 ;
        RECT 118.300 144.500 121.000 144.800 ;
        RECT 118.300 144.400 118.700 144.500 ;
        RECT 120.600 144.400 121.000 144.500 ;
        RECT 117.500 143.700 117.900 143.800 ;
        RECT 118.900 143.700 119.300 143.800 ;
        RECT 115.800 143.100 116.200 143.500 ;
        RECT 117.500 143.400 119.300 143.700 ;
        RECT 117.900 143.100 118.200 143.400 ;
        RECT 120.600 143.100 121.000 143.500 ;
        RECT 115.500 141.100 116.100 143.100 ;
        RECT 117.800 141.100 118.200 143.100 ;
        RECT 120.000 142.800 121.000 143.100 ;
        RECT 120.000 141.100 120.400 142.800 ;
        RECT 122.200 141.100 122.600 145.300 ;
        RECT 123.800 145.100 124.100 146.800 ;
        RECT 125.400 145.800 125.800 147.200 ;
        RECT 127.100 146.900 127.500 147.200 ;
        RECT 128.700 146.900 129.100 147.200 ;
        RECT 130.500 146.900 130.900 147.200 ;
        RECT 126.200 146.500 127.500 146.900 ;
        RECT 127.900 146.500 129.100 146.900 ;
        RECT 129.600 146.500 130.900 146.900 ;
        RECT 127.100 145.800 127.500 146.500 ;
        RECT 128.700 145.800 129.100 146.500 ;
        RECT 130.500 145.800 130.900 146.500 ;
        RECT 125.400 145.400 126.600 145.800 ;
        RECT 127.100 145.400 128.200 145.800 ;
        RECT 128.700 145.400 129.800 145.800 ;
        RECT 130.500 145.400 131.400 145.800 ;
        RECT 123.300 144.700 124.200 145.100 ;
        RECT 123.300 141.100 123.700 144.700 ;
        RECT 126.200 141.100 126.600 145.400 ;
        RECT 127.800 141.100 128.200 145.400 ;
        RECT 129.400 141.100 129.800 145.400 ;
        RECT 131.000 141.100 131.400 145.400 ;
        RECT 132.600 145.700 133.000 147.400 ;
        RECT 136.100 147.100 136.500 147.200 ;
        RECT 139.000 147.100 139.300 148.200 ;
        RECT 141.400 147.500 141.800 149.900 ;
        RECT 143.000 147.600 143.400 149.900 ;
        RECT 144.600 147.600 145.000 149.900 ;
        RECT 146.200 147.600 146.600 149.900 ;
        RECT 147.800 147.600 148.200 149.900 ;
        RECT 143.000 147.200 143.900 147.600 ;
        RECT 144.600 147.200 145.700 147.600 ;
        RECT 146.200 147.200 147.300 147.600 ;
        RECT 147.800 147.200 149.000 147.600 ;
        RECT 151.000 147.500 151.400 149.900 ;
        RECT 153.200 149.200 153.600 149.900 ;
        RECT 152.600 148.900 153.600 149.200 ;
        RECT 155.400 148.900 155.800 149.900 ;
        RECT 157.500 149.200 158.100 149.900 ;
        RECT 157.400 148.900 158.100 149.200 ;
        RECT 152.600 148.500 153.000 148.900 ;
        RECT 155.400 148.600 155.700 148.900 ;
        RECT 153.400 148.200 153.800 148.600 ;
        RECT 154.300 148.300 155.700 148.600 ;
        RECT 157.400 148.500 157.800 148.900 ;
        RECT 154.300 148.200 154.700 148.300 ;
        RECT 140.600 147.100 141.400 147.200 ;
        RECT 135.900 146.800 141.400 147.100 ;
        RECT 143.500 146.900 143.900 147.200 ;
        RECT 145.300 146.900 145.700 147.200 ;
        RECT 146.900 146.900 147.300 147.200 ;
        RECT 135.000 146.400 135.400 146.500 ;
        RECT 133.500 146.100 135.400 146.400 ;
        RECT 135.900 146.200 136.200 146.800 ;
        RECT 139.500 146.700 139.900 146.800 ;
        RECT 143.500 146.500 144.800 146.900 ;
        RECT 145.300 146.500 146.500 146.900 ;
        RECT 146.900 146.500 148.200 146.900 ;
        RECT 139.000 146.200 139.400 146.300 ;
        RECT 140.300 146.200 140.700 146.300 ;
        RECT 133.500 146.000 133.900 146.100 ;
        RECT 135.800 145.800 136.200 146.200 ;
        RECT 138.200 145.900 140.700 146.200 ;
        RECT 138.200 145.800 138.600 145.900 ;
        RECT 143.500 145.800 143.900 146.500 ;
        RECT 145.300 145.800 145.700 146.500 ;
        RECT 146.900 145.800 147.300 146.500 ;
        RECT 148.600 145.800 149.000 147.200 ;
        RECT 151.400 147.100 152.200 147.200 ;
        RECT 153.500 147.100 153.800 148.200 ;
        RECT 158.300 147.700 158.700 147.800 ;
        RECT 159.800 147.700 160.200 149.900 ;
        RECT 161.900 149.200 162.300 149.900 ;
        RECT 161.900 148.800 162.600 149.200 ;
        RECT 161.900 148.200 162.300 148.800 ;
        RECT 158.300 147.400 160.200 147.700 ;
        RECT 161.400 147.900 162.300 148.200 ;
        RECT 163.000 148.500 163.400 149.500 ;
        RECT 156.300 147.100 156.700 147.200 ;
        RECT 151.400 146.800 156.900 147.100 ;
        RECT 152.900 146.700 153.300 146.800 ;
        RECT 152.100 146.200 152.500 146.300 ;
        RECT 152.100 145.900 154.600 146.200 ;
        RECT 154.200 145.800 154.600 145.900 ;
        RECT 134.300 145.700 134.700 145.800 ;
        RECT 132.600 145.400 134.700 145.700 ;
        RECT 132.600 141.100 133.000 145.400 ;
        RECT 135.900 145.200 136.200 145.800 ;
        RECT 139.000 145.500 141.800 145.600 ;
        RECT 138.900 145.400 141.800 145.500 ;
        RECT 135.000 144.900 136.200 145.200 ;
        RECT 136.900 145.300 141.800 145.400 ;
        RECT 136.900 145.100 139.300 145.300 ;
        RECT 135.000 144.400 135.300 144.900 ;
        RECT 134.600 144.000 135.300 144.400 ;
        RECT 136.100 144.500 136.500 144.600 ;
        RECT 136.900 144.500 137.200 145.100 ;
        RECT 136.100 144.200 137.200 144.500 ;
        RECT 137.500 144.500 140.200 144.800 ;
        RECT 137.500 144.400 137.900 144.500 ;
        RECT 139.800 144.400 140.200 144.500 ;
        RECT 136.700 143.700 137.100 143.800 ;
        RECT 138.100 143.700 138.500 143.800 ;
        RECT 135.000 143.100 135.400 143.500 ;
        RECT 136.700 143.400 138.500 143.700 ;
        RECT 137.100 143.100 137.400 143.400 ;
        RECT 139.800 143.100 140.200 143.500 ;
        RECT 134.700 141.100 135.300 143.100 ;
        RECT 137.000 141.100 137.400 143.100 ;
        RECT 139.200 142.800 140.200 143.100 ;
        RECT 139.200 141.100 139.600 142.800 ;
        RECT 141.400 141.100 141.800 145.300 ;
        RECT 143.000 145.400 143.900 145.800 ;
        RECT 144.600 145.400 145.700 145.800 ;
        RECT 146.200 145.400 147.300 145.800 ;
        RECT 147.800 145.400 149.000 145.800 ;
        RECT 151.000 145.500 153.800 145.600 ;
        RECT 151.000 145.400 153.900 145.500 ;
        RECT 143.000 141.100 143.400 145.400 ;
        RECT 144.600 141.100 145.000 145.400 ;
        RECT 146.200 141.100 146.600 145.400 ;
        RECT 147.800 141.100 148.200 145.400 ;
        RECT 151.000 145.300 155.900 145.400 ;
        RECT 151.000 141.100 151.400 145.300 ;
        RECT 153.500 145.100 155.900 145.300 ;
        RECT 152.600 144.500 155.300 144.800 ;
        RECT 152.600 144.400 153.000 144.500 ;
        RECT 154.900 144.400 155.300 144.500 ;
        RECT 155.600 144.500 155.900 145.100 ;
        RECT 156.600 145.200 156.900 146.800 ;
        RECT 157.400 146.400 157.800 146.500 ;
        RECT 157.400 146.100 159.300 146.400 ;
        RECT 158.900 146.000 159.300 146.100 ;
        RECT 158.100 145.700 158.500 145.800 ;
        RECT 159.800 145.700 160.200 147.400 ;
        RECT 160.600 146.800 161.000 147.600 ;
        RECT 158.100 145.400 160.200 145.700 ;
        RECT 156.600 144.900 157.800 145.200 ;
        RECT 156.300 144.500 156.700 144.600 ;
        RECT 155.600 144.200 156.700 144.500 ;
        RECT 157.500 144.400 157.800 144.900 ;
        RECT 157.500 144.000 158.200 144.400 ;
        RECT 154.300 143.700 154.700 143.800 ;
        RECT 155.700 143.700 156.100 143.800 ;
        RECT 152.600 143.100 153.000 143.500 ;
        RECT 154.300 143.400 156.100 143.700 ;
        RECT 155.400 143.100 155.700 143.400 ;
        RECT 157.400 143.100 157.800 143.500 ;
        RECT 152.600 142.800 153.600 143.100 ;
        RECT 153.200 141.100 153.600 142.800 ;
        RECT 155.400 141.100 155.800 143.100 ;
        RECT 157.500 141.100 158.100 143.100 ;
        RECT 159.800 141.100 160.200 145.400 ;
        RECT 161.400 141.100 161.800 147.900 ;
        RECT 163.000 147.400 163.300 148.500 ;
        RECT 165.100 148.000 165.500 149.500 ;
        RECT 168.600 148.900 169.000 149.900 ;
        RECT 171.000 148.900 171.400 149.900 ;
        RECT 165.100 147.700 165.900 148.000 ;
        RECT 165.500 147.500 165.900 147.700 ;
        RECT 163.000 147.100 165.100 147.400 ;
        RECT 164.600 146.900 165.100 147.100 ;
        RECT 165.600 147.200 165.900 147.500 ;
        RECT 168.600 147.200 168.900 148.900 ;
        RECT 171.000 147.200 171.300 148.900 ;
        RECT 171.800 147.800 172.200 148.600 ;
        RECT 172.600 147.500 173.000 149.900 ;
        RECT 174.800 149.200 175.200 149.900 ;
        RECT 174.200 148.900 175.200 149.200 ;
        RECT 177.000 148.900 177.400 149.900 ;
        RECT 179.100 149.200 179.700 149.900 ;
        RECT 179.000 148.900 179.700 149.200 ;
        RECT 174.200 148.500 174.600 148.900 ;
        RECT 177.000 148.600 177.300 148.900 ;
        RECT 175.000 147.800 175.400 148.600 ;
        RECT 175.900 148.300 177.300 148.600 ;
        RECT 179.000 148.500 179.400 148.900 ;
        RECT 175.900 148.200 176.300 148.300 ;
        RECT 163.000 145.800 163.400 146.600 ;
        RECT 163.800 145.800 164.200 146.600 ;
        RECT 164.600 146.500 165.300 146.900 ;
        RECT 165.600 146.800 166.600 147.200 ;
        RECT 167.000 147.100 167.400 147.200 ;
        RECT 168.600 147.100 169.000 147.200 ;
        RECT 167.000 146.800 169.000 147.100 ;
        RECT 171.000 146.800 171.400 147.200 ;
        RECT 173.000 147.100 173.800 147.200 ;
        RECT 175.100 147.100 175.400 147.800 ;
        RECT 179.900 147.700 180.300 147.800 ;
        RECT 181.400 147.700 181.800 149.900 ;
        RECT 179.900 147.400 181.800 147.700 ;
        RECT 182.200 147.500 182.600 149.900 ;
        RECT 184.400 149.200 184.800 149.900 ;
        RECT 183.800 148.900 184.800 149.200 ;
        RECT 186.600 148.900 187.000 149.900 ;
        RECT 188.700 149.200 189.300 149.900 ;
        RECT 188.600 148.900 189.300 149.200 ;
        RECT 183.800 148.500 184.200 148.900 ;
        RECT 186.600 148.600 186.900 148.900 ;
        RECT 184.600 148.200 185.000 148.600 ;
        RECT 185.500 148.300 186.900 148.600 ;
        RECT 188.600 148.500 189.000 148.900 ;
        RECT 185.500 148.200 185.900 148.300 ;
        RECT 175.800 147.100 176.200 147.200 ;
        RECT 177.900 147.100 178.300 147.200 ;
        RECT 173.000 146.800 178.500 147.100 ;
        RECT 164.600 145.500 164.900 146.500 ;
        RECT 163.000 145.200 164.900 145.500 ;
        RECT 165.600 145.200 165.900 146.800 ;
        RECT 162.200 144.400 162.600 145.200 ;
        RECT 163.000 143.500 163.300 145.200 ;
        RECT 165.400 144.900 165.900 145.200 ;
        RECT 168.600 145.100 168.900 146.800 ;
        RECT 170.200 145.400 170.600 146.200 ;
        RECT 171.000 145.200 171.300 146.800 ;
        RECT 174.500 146.700 174.900 146.800 ;
        RECT 173.700 146.200 174.100 146.300 ;
        RECT 175.000 146.200 175.400 146.300 ;
        RECT 173.700 145.900 176.200 146.200 ;
        RECT 175.800 145.800 176.200 145.900 ;
        RECT 172.600 145.500 175.400 145.600 ;
        RECT 172.600 145.400 175.500 145.500 ;
        RECT 172.600 145.300 177.500 145.400 ;
        RECT 171.000 145.100 171.400 145.200 ;
        RECT 165.100 144.600 165.900 144.900 ;
        RECT 168.100 144.700 169.000 145.100 ;
        RECT 170.500 144.700 171.400 145.100 ;
        RECT 163.000 141.500 163.400 143.500 ;
        RECT 165.100 141.100 165.500 144.600 ;
        RECT 168.100 141.100 168.500 144.700 ;
        RECT 170.500 141.100 170.900 144.700 ;
        RECT 172.600 141.100 173.000 145.300 ;
        RECT 175.100 145.100 177.500 145.300 ;
        RECT 174.200 144.500 176.900 144.800 ;
        RECT 174.200 144.400 174.600 144.500 ;
        RECT 176.500 144.400 176.900 144.500 ;
        RECT 177.200 144.500 177.500 145.100 ;
        RECT 178.200 145.200 178.500 146.800 ;
        RECT 179.000 146.400 179.400 146.500 ;
        RECT 179.000 146.100 180.900 146.400 ;
        RECT 180.500 146.000 180.900 146.100 ;
        RECT 179.700 145.700 180.100 145.800 ;
        RECT 181.400 145.700 181.800 147.400 ;
        RECT 182.600 147.100 183.400 147.200 ;
        RECT 184.700 147.100 185.000 148.200 ;
        RECT 189.500 147.700 189.900 147.800 ;
        RECT 191.000 147.700 191.400 149.900 ;
        RECT 189.500 147.400 191.400 147.700 ;
        RECT 187.500 147.100 187.900 147.200 ;
        RECT 182.600 146.800 188.100 147.100 ;
        RECT 184.100 146.700 184.500 146.800 ;
        RECT 183.300 146.200 183.700 146.300 ;
        RECT 184.600 146.200 185.000 146.300 ;
        RECT 183.300 145.900 185.800 146.200 ;
        RECT 185.400 145.800 185.800 145.900 ;
        RECT 179.700 145.400 181.800 145.700 ;
        RECT 178.200 144.900 179.400 145.200 ;
        RECT 177.900 144.500 178.300 144.600 ;
        RECT 177.200 144.200 178.300 144.500 ;
        RECT 179.100 144.400 179.400 144.900 ;
        RECT 179.100 144.000 179.800 144.400 ;
        RECT 175.900 143.700 176.300 143.800 ;
        RECT 177.300 143.700 177.700 143.800 ;
        RECT 174.200 143.100 174.600 143.500 ;
        RECT 175.900 143.400 177.700 143.700 ;
        RECT 177.000 143.100 177.300 143.400 ;
        RECT 179.000 143.100 179.400 143.500 ;
        RECT 174.200 142.800 175.200 143.100 ;
        RECT 174.800 141.100 175.200 142.800 ;
        RECT 177.000 141.100 177.400 143.100 ;
        RECT 179.100 141.100 179.700 143.100 ;
        RECT 181.400 141.100 181.800 145.400 ;
        RECT 182.200 145.500 185.000 145.600 ;
        RECT 182.200 145.400 185.100 145.500 ;
        RECT 182.200 145.300 187.100 145.400 ;
        RECT 182.200 141.100 182.600 145.300 ;
        RECT 184.700 145.100 187.100 145.300 ;
        RECT 183.800 144.500 186.500 144.800 ;
        RECT 183.800 144.400 184.200 144.500 ;
        RECT 186.100 144.400 186.500 144.500 ;
        RECT 186.800 144.500 187.100 145.100 ;
        RECT 187.800 145.200 188.100 146.800 ;
        RECT 188.600 146.400 189.000 146.500 ;
        RECT 188.600 146.100 190.500 146.400 ;
        RECT 190.100 146.000 190.500 146.100 ;
        RECT 189.300 145.700 189.700 145.800 ;
        RECT 191.000 145.700 191.400 147.400 ;
        RECT 191.800 147.600 192.200 149.900 ;
        RECT 191.800 147.300 192.900 147.600 ;
        RECT 189.300 145.400 191.400 145.700 ;
        RECT 187.800 144.900 189.000 145.200 ;
        RECT 187.500 144.500 187.900 144.600 ;
        RECT 186.800 144.200 187.900 144.500 ;
        RECT 188.700 144.400 189.000 144.900 ;
        RECT 188.700 144.000 189.400 144.400 ;
        RECT 185.500 143.700 185.900 143.800 ;
        RECT 186.900 143.700 187.300 143.800 ;
        RECT 183.800 143.100 184.200 143.500 ;
        RECT 185.500 143.400 187.300 143.700 ;
        RECT 186.600 143.100 186.900 143.400 ;
        RECT 188.600 143.100 189.000 143.500 ;
        RECT 183.800 142.800 184.800 143.100 ;
        RECT 184.400 141.100 184.800 142.800 ;
        RECT 186.600 141.100 187.000 143.100 ;
        RECT 188.700 141.100 189.300 143.100 ;
        RECT 191.000 141.100 191.400 145.400 ;
        RECT 192.600 145.800 192.900 147.300 ;
        RECT 193.400 146.200 193.800 149.900 ;
        RECT 192.600 145.400 193.200 145.800 ;
        RECT 192.600 145.100 192.900 145.400 ;
        RECT 193.500 145.100 193.800 146.200 ;
        RECT 191.800 144.800 192.900 145.100 ;
        RECT 191.800 141.100 192.200 144.800 ;
        RECT 193.400 141.100 193.800 145.100 ;
        RECT 0.600 135.600 1.000 139.900 ;
        RECT 2.700 137.900 3.300 139.900 ;
        RECT 5.000 137.900 5.400 139.900 ;
        RECT 7.200 138.200 7.600 139.900 ;
        RECT 7.200 137.900 8.200 138.200 ;
        RECT 3.000 137.500 3.400 137.900 ;
        RECT 5.100 137.600 5.400 137.900 ;
        RECT 4.700 137.300 6.500 137.600 ;
        RECT 7.800 137.500 8.200 137.900 ;
        RECT 4.700 137.200 5.100 137.300 ;
        RECT 6.100 137.200 6.500 137.300 ;
        RECT 2.600 136.600 3.300 137.000 ;
        RECT 3.000 136.100 3.300 136.600 ;
        RECT 4.100 136.500 5.200 136.800 ;
        RECT 4.100 136.400 4.500 136.500 ;
        RECT 3.000 135.800 4.200 136.100 ;
        RECT 0.600 135.300 2.700 135.600 ;
        RECT 0.600 133.600 1.000 135.300 ;
        RECT 2.300 135.200 2.700 135.300 ;
        RECT 1.500 134.900 1.900 135.000 ;
        RECT 1.500 134.600 3.400 134.900 ;
        RECT 3.000 134.500 3.400 134.600 ;
        RECT 3.900 134.200 4.200 135.800 ;
        RECT 4.900 135.900 5.200 136.500 ;
        RECT 5.500 136.500 5.900 136.600 ;
        RECT 7.800 136.500 8.200 136.600 ;
        RECT 5.500 136.200 8.200 136.500 ;
        RECT 4.900 135.700 7.300 135.900 ;
        RECT 9.400 135.700 9.800 139.900 ;
        RECT 4.900 135.600 9.800 135.700 ;
        RECT 6.900 135.500 9.800 135.600 ;
        RECT 7.000 135.400 9.800 135.500 ;
        RECT 10.200 135.700 10.600 139.900 ;
        RECT 12.400 138.200 12.800 139.900 ;
        RECT 11.800 137.900 12.800 138.200 ;
        RECT 14.600 137.900 15.000 139.900 ;
        RECT 16.700 137.900 17.300 139.900 ;
        RECT 11.800 137.500 12.200 137.900 ;
        RECT 14.600 137.600 14.900 137.900 ;
        RECT 13.500 137.300 15.300 137.600 ;
        RECT 16.600 137.500 17.000 137.900 ;
        RECT 13.500 137.200 13.900 137.300 ;
        RECT 14.900 137.200 15.300 137.300 ;
        RECT 11.800 136.500 12.200 136.600 ;
        RECT 14.100 136.500 14.500 136.600 ;
        RECT 11.800 136.200 14.500 136.500 ;
        RECT 14.800 136.500 15.900 136.800 ;
        RECT 14.800 135.900 15.100 136.500 ;
        RECT 15.500 136.400 15.900 136.500 ;
        RECT 16.700 136.600 17.400 137.000 ;
        RECT 16.700 136.100 17.000 136.600 ;
        RECT 12.700 135.700 15.100 135.900 ;
        RECT 10.200 135.600 15.100 135.700 ;
        RECT 15.800 135.800 17.000 136.100 ;
        RECT 10.200 135.500 13.100 135.600 ;
        RECT 10.200 135.400 13.000 135.500 ;
        RECT 6.200 135.100 6.600 135.200 ;
        RECT 13.400 135.100 13.800 135.200 ;
        RECT 6.200 134.800 8.700 135.100 ;
        RECT 8.300 134.700 8.700 134.800 ;
        RECT 11.300 134.800 13.800 135.100 ;
        RECT 11.300 134.700 11.700 134.800 ;
        RECT 7.500 134.200 7.900 134.300 ;
        RECT 12.100 134.200 12.500 134.300 ;
        RECT 15.800 134.200 16.100 135.800 ;
        RECT 19.000 135.600 19.400 139.900 ;
        RECT 21.100 136.300 21.500 139.900 ;
        RECT 20.600 135.900 21.500 136.300 ;
        RECT 22.200 137.500 22.600 139.500 ;
        RECT 17.300 135.300 19.400 135.600 ;
        RECT 17.300 135.200 17.700 135.300 ;
        RECT 18.100 134.900 18.500 135.000 ;
        RECT 16.600 134.600 18.500 134.900 ;
        RECT 16.600 134.500 17.000 134.600 ;
        RECT 3.900 133.900 9.400 134.200 ;
        RECT 4.100 133.800 4.500 133.900 ;
        RECT 7.000 133.800 7.400 133.900 ;
        RECT 8.600 133.800 9.400 133.900 ;
        RECT 10.600 133.900 16.100 134.200 ;
        RECT 10.600 133.800 11.400 133.900 ;
        RECT 0.600 133.300 2.500 133.600 ;
        RECT 0.600 131.100 1.000 133.300 ;
        RECT 2.100 133.200 2.500 133.300 ;
        RECT 7.000 132.800 7.300 133.800 ;
        RECT 6.100 132.700 6.500 132.800 ;
        RECT 3.000 132.100 3.400 132.500 ;
        RECT 5.100 132.400 6.500 132.700 ;
        RECT 7.000 132.400 7.400 132.800 ;
        RECT 5.100 132.100 5.400 132.400 ;
        RECT 7.800 132.100 8.200 132.500 ;
        RECT 2.700 131.800 3.400 132.100 ;
        RECT 2.700 131.100 3.300 131.800 ;
        RECT 5.000 131.100 5.400 132.100 ;
        RECT 7.200 131.800 8.200 132.100 ;
        RECT 7.200 131.100 7.600 131.800 ;
        RECT 9.400 131.100 9.800 133.500 ;
        RECT 10.200 131.100 10.600 133.500 ;
        RECT 12.700 132.800 13.000 133.900 ;
        RECT 14.200 133.800 14.600 133.900 ;
        RECT 15.500 133.800 15.900 133.900 ;
        RECT 19.000 133.600 19.400 135.300 ;
        RECT 19.800 134.800 20.200 135.200 ;
        RECT 19.800 134.100 20.100 134.800 ;
        RECT 20.700 134.200 21.000 135.900 ;
        RECT 22.200 135.800 22.500 137.500 ;
        RECT 24.300 136.400 24.700 139.900 ;
        RECT 24.300 136.100 25.100 136.400 ;
        RECT 21.400 134.800 21.800 135.600 ;
        RECT 22.200 135.500 24.100 135.800 ;
        RECT 22.200 134.400 22.600 135.200 ;
        RECT 23.000 134.400 23.400 135.200 ;
        RECT 23.800 134.500 24.100 135.500 ;
        RECT 20.600 134.100 21.000 134.200 ;
        RECT 19.800 133.800 21.000 134.100 ;
        RECT 23.800 134.100 24.500 134.500 ;
        RECT 24.800 134.200 25.100 136.100 ;
        RECT 27.000 136.200 27.400 139.900 ;
        RECT 27.000 135.900 28.100 136.200 ;
        RECT 28.600 135.900 29.000 139.900 ;
        RECT 29.700 136.300 30.100 139.900 ;
        RECT 33.700 136.400 34.100 139.900 ;
        RECT 35.800 137.500 36.200 139.500 ;
        RECT 29.700 135.900 30.600 136.300 ;
        RECT 33.300 136.100 34.100 136.400 ;
        RECT 27.800 135.600 28.100 135.900 ;
        RECT 25.400 135.100 25.800 135.600 ;
        RECT 27.800 135.200 28.400 135.600 ;
        RECT 26.200 135.100 26.600 135.200 ;
        RECT 25.400 134.800 26.600 135.100 ;
        RECT 23.800 133.900 24.300 134.100 ;
        RECT 17.500 133.300 19.400 133.600 ;
        RECT 17.500 133.200 17.900 133.300 ;
        RECT 11.800 132.100 12.200 132.500 ;
        RECT 12.600 132.400 13.000 132.800 ;
        RECT 13.500 132.700 13.900 132.800 ;
        RECT 13.500 132.400 14.900 132.700 ;
        RECT 14.600 132.100 14.900 132.400 ;
        RECT 16.600 132.100 17.000 132.500 ;
        RECT 11.800 131.800 12.800 132.100 ;
        RECT 12.400 131.100 12.800 131.800 ;
        RECT 14.600 131.100 15.000 132.100 ;
        RECT 16.600 131.800 17.300 132.100 ;
        RECT 16.700 131.100 17.300 131.800 ;
        RECT 19.000 131.100 19.400 133.300 ;
        RECT 19.800 132.400 20.200 133.200 ;
        RECT 20.700 132.100 21.000 133.800 ;
        RECT 20.600 131.100 21.000 132.100 ;
        RECT 22.200 133.600 24.300 133.900 ;
        RECT 24.800 133.800 25.800 134.200 ;
        RECT 22.200 132.500 22.500 133.600 ;
        RECT 24.800 133.500 25.100 133.800 ;
        RECT 27.800 133.700 28.100 135.200 ;
        RECT 28.700 134.800 29.000 135.900 ;
        RECT 29.400 134.800 29.800 135.600 ;
        RECT 24.700 133.300 25.100 133.500 ;
        RECT 24.300 133.200 25.100 133.300 ;
        RECT 23.800 133.000 25.100 133.200 ;
        RECT 27.000 133.400 28.100 133.700 ;
        RECT 23.800 132.800 24.700 133.000 ;
        RECT 22.200 131.500 22.600 132.500 ;
        RECT 24.300 131.500 24.700 132.800 ;
        RECT 27.000 131.100 27.400 133.400 ;
        RECT 28.600 131.100 29.000 134.800 ;
        RECT 30.200 134.200 30.500 135.900 ;
        RECT 32.600 134.800 33.000 135.600 ;
        RECT 33.300 134.200 33.600 136.100 ;
        RECT 35.900 135.800 36.200 137.500 ;
        RECT 37.000 136.800 37.400 137.200 ;
        RECT 37.000 136.200 37.300 136.800 ;
        RECT 37.700 136.200 38.100 139.900 ;
        RECT 36.600 135.900 37.300 136.200 ;
        RECT 37.600 135.900 38.100 136.200 ;
        RECT 39.800 135.900 40.200 139.900 ;
        RECT 40.600 136.200 41.000 139.900 ;
        RECT 42.200 136.200 42.600 139.900 ;
        RECT 43.800 137.900 44.200 139.900 ;
        RECT 43.900 137.800 44.200 137.900 ;
        RECT 45.400 137.900 45.800 139.900 ;
        RECT 45.400 137.800 45.700 137.900 ;
        RECT 43.900 137.500 45.700 137.800 ;
        RECT 44.600 136.400 45.000 137.200 ;
        RECT 45.400 136.200 45.700 137.500 ;
        RECT 47.800 136.200 48.200 139.900 ;
        RECT 50.000 139.200 50.800 139.900 ;
        RECT 50.000 138.800 51.400 139.200 ;
        RECT 48.600 136.200 49.000 136.300 ;
        RECT 50.000 136.200 50.800 138.800 ;
        RECT 40.600 135.900 42.600 136.200 ;
        RECT 36.600 135.800 37.000 135.900 ;
        RECT 34.300 135.500 36.200 135.800 ;
        RECT 34.300 134.500 34.600 135.500 ;
        RECT 30.200 133.800 30.600 134.200 ;
        RECT 31.800 134.100 32.200 134.200 ;
        RECT 32.600 134.100 33.600 134.200 ;
        RECT 33.900 134.100 34.600 134.500 ;
        RECT 35.000 134.400 35.400 135.200 ;
        RECT 35.800 134.400 36.200 135.200 ;
        RECT 37.600 134.200 37.900 135.900 ;
        RECT 39.900 135.200 40.200 135.900 ;
        RECT 43.000 135.400 43.400 136.200 ;
        RECT 45.400 135.800 45.800 136.200 ;
        RECT 47.800 135.900 49.000 136.200 ;
        RECT 49.800 135.900 50.800 136.200 ;
        RECT 51.900 136.200 52.300 136.300 ;
        RECT 52.600 136.200 53.000 139.900 ;
        RECT 54.200 136.400 54.600 139.900 ;
        RECT 51.900 135.900 53.000 136.200 ;
        RECT 54.100 135.900 54.600 136.400 ;
        RECT 55.800 136.200 56.200 139.900 ;
        RECT 54.900 135.900 56.200 136.200 ;
        RECT 57.900 136.200 58.300 139.900 ;
        RECT 60.900 139.200 61.300 139.900 ;
        RECT 60.900 138.800 61.800 139.200 ;
        RECT 58.600 136.800 59.000 137.200 ;
        RECT 58.700 136.200 59.000 136.800 ;
        RECT 60.200 136.800 60.600 137.200 ;
        RECT 60.200 136.200 60.500 136.800 ;
        RECT 60.900 136.200 61.300 138.800 ;
        RECT 63.800 137.800 64.200 139.900 ;
        RECT 65.400 137.900 65.800 139.900 ;
        RECT 67.000 137.900 67.400 139.900 ;
        RECT 65.400 137.800 65.700 137.900 ;
        RECT 63.900 137.500 65.700 137.800 ;
        RECT 67.100 137.800 67.400 137.900 ;
        RECT 68.600 137.900 69.000 139.900 ;
        RECT 68.600 137.800 68.900 137.900 ;
        RECT 67.100 137.500 68.900 137.800 ;
        RECT 64.600 136.400 65.000 137.200 ;
        RECT 65.400 136.200 65.700 137.500 ;
        RECT 67.800 136.400 68.200 137.200 ;
        RECT 68.600 136.200 68.900 137.500 ;
        RECT 57.900 135.900 58.400 136.200 ;
        RECT 58.700 135.900 59.400 136.200 ;
        RECT 41.800 135.200 42.200 135.400 ;
        RECT 38.200 134.400 38.600 135.200 ;
        RECT 39.800 134.900 41.000 135.200 ;
        RECT 41.800 134.900 42.600 135.200 ;
        RECT 39.800 134.800 40.200 134.900 ;
        RECT 31.800 133.800 33.600 134.100 ;
        RECT 30.200 132.200 30.500 133.800 ;
        RECT 33.300 133.500 33.600 133.800 ;
        RECT 34.100 133.900 34.600 134.100 ;
        RECT 34.100 133.600 36.200 133.900 ;
        RECT 36.600 133.800 37.900 134.200 ;
        RECT 39.000 134.100 39.400 134.200 ;
        RECT 38.600 133.800 39.400 134.100 ;
        RECT 33.300 133.300 33.700 133.500 ;
        RECT 31.000 132.400 31.400 133.200 ;
        RECT 33.300 133.000 34.100 133.300 ;
        RECT 30.200 131.100 30.600 132.200 ;
        RECT 33.700 131.500 34.100 133.000 ;
        RECT 35.900 132.500 36.200 133.600 ;
        RECT 36.700 133.100 37.000 133.800 ;
        RECT 38.600 133.600 39.000 133.800 ;
        RECT 37.500 133.100 39.300 133.300 ;
        RECT 35.800 131.500 36.200 132.500 ;
        RECT 36.600 131.100 37.000 133.100 ;
        RECT 37.400 133.000 39.400 133.100 ;
        RECT 37.400 131.100 37.800 133.000 ;
        RECT 39.000 131.100 39.400 133.000 ;
        RECT 39.800 132.800 40.200 133.200 ;
        RECT 40.700 133.100 41.000 134.900 ;
        RECT 42.200 134.800 42.600 134.900 ;
        RECT 43.800 134.800 45.000 135.200 ;
        RECT 41.400 133.800 41.800 134.600 ;
        RECT 45.400 134.200 45.700 135.800 ;
        RECT 49.800 135.200 50.100 135.900 ;
        RECT 51.900 135.600 52.200 135.900 ;
        RECT 50.500 135.300 52.200 135.600 ;
        RECT 50.500 135.200 50.900 135.300 ;
        RECT 49.400 134.900 50.100 135.200 ;
        RECT 51.600 134.900 52.000 135.000 ;
        RECT 49.400 134.800 50.300 134.900 ;
        RECT 49.800 134.600 50.300 134.800 ;
        RECT 44.900 134.100 45.700 134.200 ;
        RECT 43.800 133.900 45.700 134.100 ;
        RECT 43.800 133.800 45.200 133.900 ;
        RECT 47.800 133.800 48.600 134.200 ;
        RECT 49.200 133.800 49.600 134.200 ;
        RECT 39.900 132.400 40.300 132.800 ;
        RECT 40.600 131.100 41.000 133.100 ;
        RECT 43.800 133.200 44.100 133.800 ;
        RECT 43.800 132.800 44.200 133.200 ;
        RECT 44.800 131.100 45.200 133.800 ;
        RECT 49.300 133.600 49.600 133.800 ;
        RECT 48.600 133.400 49.000 133.500 ;
        RECT 47.800 133.100 49.000 133.400 ;
        RECT 49.300 133.200 49.700 133.600 ;
        RECT 47.800 131.100 48.200 133.100 ;
        RECT 50.000 132.900 50.300 134.600 ;
        RECT 50.700 134.600 52.000 134.900 ;
        RECT 50.700 134.300 51.000 134.600 ;
        RECT 50.600 133.900 51.000 134.300 ;
        RECT 54.100 134.200 54.400 135.900 ;
        RECT 54.900 134.900 55.200 135.900 ;
        RECT 54.700 134.500 55.200 134.900 ;
        RECT 52.200 134.100 53.000 134.200 ;
        RECT 51.300 133.800 53.000 134.100 ;
        RECT 54.100 133.800 54.600 134.200 ;
        RECT 51.300 133.600 51.600 133.800 ;
        RECT 50.600 133.300 51.600 133.600 ;
        RECT 51.900 133.400 52.300 133.500 ;
        RECT 50.600 133.200 51.400 133.300 ;
        RECT 51.900 133.100 53.000 133.400 ;
        RECT 50.000 131.100 50.800 132.900 ;
        RECT 52.600 131.100 53.000 133.100 ;
        RECT 54.100 133.100 54.400 133.800 ;
        RECT 54.900 133.700 55.200 134.500 ;
        RECT 55.700 134.800 56.200 135.200 ;
        RECT 55.700 134.400 56.100 134.800 ;
        RECT 57.400 134.400 57.800 135.200 ;
        RECT 58.100 135.100 58.400 135.900 ;
        RECT 59.000 135.800 59.400 135.900 ;
        RECT 59.800 135.900 60.500 136.200 ;
        RECT 60.800 135.900 61.300 136.200 ;
        RECT 59.800 135.800 60.200 135.900 ;
        RECT 59.800 135.100 60.100 135.800 ;
        RECT 58.100 134.800 60.100 135.100 ;
        RECT 58.100 134.200 58.400 134.800 ;
        RECT 60.800 134.200 61.100 135.900 ;
        RECT 63.000 135.400 63.400 136.200 ;
        RECT 65.400 135.800 65.800 136.200 ;
        RECT 61.400 134.400 61.800 135.200 ;
        RECT 63.800 134.800 64.600 135.200 ;
        RECT 65.400 134.200 65.700 135.800 ;
        RECT 66.200 135.400 66.600 136.200 ;
        RECT 68.600 135.800 69.000 136.200 ;
        RECT 67.000 134.800 67.800 135.200 ;
        RECT 68.600 134.200 68.900 135.800 ;
        RECT 56.600 134.100 57.000 134.200 ;
        RECT 56.600 133.800 57.400 134.100 ;
        RECT 58.100 133.800 59.400 134.200 ;
        RECT 59.800 133.800 61.100 134.200 ;
        RECT 62.200 134.100 62.600 134.200 ;
        RECT 64.900 134.100 65.700 134.200 ;
        RECT 68.100 134.100 68.900 134.200 ;
        RECT 61.800 133.800 62.600 134.100 ;
        RECT 64.800 133.900 65.700 134.100 ;
        RECT 68.000 133.900 68.900 134.100 ;
        RECT 54.900 133.400 56.200 133.700 ;
        RECT 57.000 133.600 57.400 133.800 ;
        RECT 54.100 132.800 54.600 133.100 ;
        RECT 54.200 131.100 54.600 132.800 ;
        RECT 55.800 131.100 56.200 133.400 ;
        RECT 56.700 133.100 58.500 133.300 ;
        RECT 59.000 133.100 59.300 133.800 ;
        RECT 59.900 133.100 60.200 133.800 ;
        RECT 61.800 133.600 62.200 133.800 ;
        RECT 60.700 133.100 62.500 133.300 ;
        RECT 56.600 133.000 58.600 133.100 ;
        RECT 56.600 131.100 57.000 133.000 ;
        RECT 58.200 131.100 58.600 133.000 ;
        RECT 59.000 131.100 59.400 133.100 ;
        RECT 59.800 131.100 60.200 133.100 ;
        RECT 60.600 133.000 62.600 133.100 ;
        RECT 60.600 131.100 61.000 133.000 ;
        RECT 62.200 131.100 62.600 133.000 ;
        RECT 64.800 131.100 65.200 133.900 ;
        RECT 68.000 131.100 68.400 133.900 ;
        RECT 69.400 133.400 69.800 134.200 ;
        RECT 70.200 133.200 70.600 139.900 ;
        RECT 72.600 137.900 73.000 139.900 ;
        RECT 72.700 137.800 73.000 137.900 ;
        RECT 74.200 137.900 74.600 139.900 ;
        RECT 74.200 137.800 74.500 137.900 ;
        RECT 72.700 137.500 74.500 137.800 ;
        RECT 71.000 135.800 71.400 136.600 ;
        RECT 73.400 136.400 73.800 137.200 ;
        RECT 74.200 136.200 74.500 137.500 ;
        RECT 75.000 136.200 75.400 139.900 ;
        RECT 77.200 139.200 78.000 139.900 ;
        RECT 77.200 138.800 78.600 139.200 ;
        RECT 75.700 136.200 76.100 136.300 ;
        RECT 71.800 135.400 72.200 136.200 ;
        RECT 74.200 135.800 74.600 136.200 ;
        RECT 75.000 135.900 76.100 136.200 ;
        RECT 77.200 136.200 78.000 138.800 ;
        RECT 79.000 136.200 79.400 136.300 ;
        RECT 79.800 136.200 80.200 139.900 ;
        RECT 77.200 135.900 78.200 136.200 ;
        RECT 79.000 135.900 80.200 136.200 ;
        RECT 80.600 137.500 81.000 139.500 ;
        RECT 82.700 139.200 83.100 139.900 ;
        RECT 82.700 138.800 83.400 139.200 ;
        RECT 72.600 134.800 73.400 135.200 ;
        RECT 74.200 134.200 74.500 135.800 ;
        RECT 75.800 135.600 76.100 135.900 ;
        RECT 75.800 135.300 77.500 135.600 ;
        RECT 77.100 135.200 77.500 135.300 ;
        RECT 77.900 135.200 78.200 135.900 ;
        RECT 80.600 135.800 80.900 137.500 ;
        RECT 82.700 136.400 83.100 138.800 ;
        RECT 82.700 136.100 83.500 136.400 ;
        RECT 80.600 135.500 82.500 135.800 ;
        RECT 76.000 134.900 76.400 135.000 ;
        RECT 77.900 134.900 78.600 135.200 ;
        RECT 76.000 134.600 77.300 134.900 ;
        RECT 77.000 134.300 77.300 134.600 ;
        RECT 77.700 134.800 78.600 134.900 ;
        RECT 77.700 134.600 78.200 134.800 ;
        RECT 71.000 133.800 71.400 134.200 ;
        RECT 73.700 134.100 74.600 134.200 ;
        RECT 73.600 133.800 74.600 134.100 ;
        RECT 75.000 134.100 75.800 134.200 ;
        RECT 75.000 133.800 76.700 134.100 ;
        RECT 77.000 133.900 77.400 134.300 ;
        RECT 71.000 133.200 71.300 133.800 ;
        RECT 70.200 132.800 71.300 133.200 ;
        RECT 70.700 131.100 71.100 132.800 ;
        RECT 73.600 131.100 74.000 133.800 ;
        RECT 76.400 133.600 76.700 133.800 ;
        RECT 75.700 133.400 76.100 133.500 ;
        RECT 75.000 133.100 76.100 133.400 ;
        RECT 76.400 133.300 77.400 133.600 ;
        RECT 76.600 133.200 77.400 133.300 ;
        RECT 75.000 131.100 75.400 133.100 ;
        RECT 77.700 132.900 78.000 134.600 ;
        RECT 80.600 134.400 81.000 135.200 ;
        RECT 81.400 134.400 81.800 135.200 ;
        RECT 82.200 134.500 82.500 135.500 ;
        RECT 78.400 133.800 78.800 134.200 ;
        RECT 79.400 133.800 80.200 134.200 ;
        RECT 82.200 134.100 82.900 134.500 ;
        RECT 83.200 134.200 83.500 136.100 ;
        RECT 85.400 136.200 85.800 139.900 ;
        RECT 87.000 136.200 87.400 139.900 ;
        RECT 85.400 135.900 87.400 136.200 ;
        RECT 87.800 135.900 88.200 139.900 ;
        RECT 89.000 136.800 89.400 137.200 ;
        RECT 89.000 136.200 89.300 136.800 ;
        RECT 89.700 136.200 90.100 139.900 ;
        RECT 93.700 139.200 94.100 139.900 ;
        RECT 93.700 138.800 94.600 139.200 ;
        RECT 93.700 136.400 94.100 138.800 ;
        RECT 95.800 137.500 96.200 139.500 ;
        RECT 88.600 135.900 89.300 136.200 ;
        RECT 89.600 135.900 90.100 136.200 ;
        RECT 93.300 136.100 94.100 136.400 ;
        RECT 83.800 134.800 84.200 135.600 ;
        RECT 85.800 135.200 86.200 135.400 ;
        RECT 87.800 135.200 88.100 135.900 ;
        RECT 88.600 135.800 89.000 135.900 ;
        RECT 85.400 134.900 86.200 135.200 ;
        RECT 87.000 134.900 88.200 135.200 ;
        RECT 85.400 134.800 85.800 134.900 ;
        RECT 82.200 133.900 82.700 134.100 ;
        RECT 78.400 133.600 78.700 133.800 ;
        RECT 78.300 133.200 78.700 133.600 ;
        RECT 80.600 133.600 82.700 133.900 ;
        RECT 83.200 133.800 84.200 134.200 ;
        RECT 84.600 134.100 85.000 134.200 ;
        RECT 86.200 134.100 86.600 134.600 ;
        RECT 84.600 133.800 86.600 134.100 ;
        RECT 79.000 133.400 79.400 133.500 ;
        RECT 79.000 133.100 80.200 133.400 ;
        RECT 77.200 131.100 78.000 132.900 ;
        RECT 79.800 131.100 80.200 133.100 ;
        RECT 80.600 132.500 80.900 133.600 ;
        RECT 83.200 133.500 83.500 133.800 ;
        RECT 83.100 133.300 83.500 133.500 ;
        RECT 82.700 133.000 83.500 133.300 ;
        RECT 87.000 133.100 87.300 134.900 ;
        RECT 87.800 134.800 88.200 134.900 ;
        RECT 89.600 134.200 89.900 135.900 ;
        RECT 90.200 134.400 90.600 135.200 ;
        RECT 92.600 134.800 93.000 135.600 ;
        RECT 93.300 134.200 93.600 136.100 ;
        RECT 95.900 135.800 96.200 137.500 ;
        RECT 99.000 136.400 99.400 139.900 ;
        RECT 94.300 135.500 96.200 135.800 ;
        RECT 98.900 135.900 99.400 136.400 ;
        RECT 100.600 136.200 101.000 139.900 ;
        RECT 99.700 135.900 101.000 136.200 ;
        RECT 101.400 137.500 101.800 139.500 ;
        RECT 103.500 139.200 103.900 139.900 ;
        RECT 108.100 139.200 108.500 139.900 ;
        RECT 103.500 138.800 104.200 139.200 ;
        RECT 108.100 138.800 109.000 139.200 ;
        RECT 94.300 134.500 94.600 135.500 ;
        RECT 88.600 133.800 89.900 134.200 ;
        RECT 91.000 134.100 91.400 134.200 ;
        RECT 90.600 133.800 91.400 134.100 ;
        RECT 92.600 133.800 93.600 134.200 ;
        RECT 93.900 134.100 94.600 134.500 ;
        RECT 95.000 134.400 95.400 135.200 ;
        RECT 95.800 135.100 96.200 135.200 ;
        RECT 96.600 135.100 97.000 135.200 ;
        RECT 95.800 134.800 97.000 135.100 ;
        RECT 95.800 134.400 96.200 134.800 ;
        RECT 87.800 133.100 88.200 133.200 ;
        RECT 88.700 133.100 89.000 133.800 ;
        RECT 90.600 133.600 91.000 133.800 ;
        RECT 93.300 133.500 93.600 133.800 ;
        RECT 94.100 133.900 94.600 134.100 ;
        RECT 96.600 134.100 96.900 134.800 ;
        RECT 98.900 134.200 99.200 135.900 ;
        RECT 99.700 134.900 100.000 135.900 ;
        RECT 101.400 135.800 101.700 137.500 ;
        RECT 103.500 136.400 103.900 138.800 ;
        RECT 108.100 136.400 108.500 138.800 ;
        RECT 110.200 137.500 110.600 139.500 ;
        RECT 103.500 136.100 104.300 136.400 ;
        RECT 101.400 135.500 103.300 135.800 ;
        RECT 99.500 134.500 100.000 134.900 ;
        RECT 98.900 134.100 99.400 134.200 ;
        RECT 94.100 133.600 96.200 133.900 ;
        RECT 96.600 133.800 99.400 134.100 ;
        RECT 93.300 133.300 93.700 133.500 ;
        RECT 89.500 133.100 91.300 133.300 ;
        RECT 80.600 131.500 81.000 132.500 ;
        RECT 82.700 131.500 83.100 133.000 ;
        RECT 87.000 131.100 87.400 133.100 ;
        RECT 87.800 132.800 89.000 133.100 ;
        RECT 87.700 132.400 88.100 132.800 ;
        RECT 88.600 131.100 89.000 132.800 ;
        RECT 89.400 133.000 91.400 133.100 ;
        RECT 93.300 133.000 94.100 133.300 ;
        RECT 89.400 131.100 89.800 133.000 ;
        RECT 91.000 131.100 91.400 133.000 ;
        RECT 93.700 131.500 94.100 133.000 ;
        RECT 95.900 132.500 96.200 133.600 ;
        RECT 98.900 133.100 99.200 133.800 ;
        RECT 99.700 133.700 100.000 134.500 ;
        RECT 100.500 134.800 101.000 135.200 ;
        RECT 100.500 134.400 100.900 134.800 ;
        RECT 101.400 134.400 101.800 135.200 ;
        RECT 102.200 134.400 102.600 135.200 ;
        RECT 103.000 134.500 103.300 135.500 ;
        RECT 103.000 134.100 103.700 134.500 ;
        RECT 104.000 134.200 104.300 136.100 ;
        RECT 107.700 136.100 108.500 136.400 ;
        RECT 104.600 134.800 105.000 135.600 ;
        RECT 107.000 134.800 107.400 135.600 ;
        RECT 107.700 134.200 108.000 136.100 ;
        RECT 110.300 135.800 110.600 137.500 ;
        RECT 108.700 135.500 110.600 135.800 ;
        RECT 108.700 134.500 109.000 135.500 ;
        RECT 103.000 133.900 103.500 134.100 ;
        RECT 99.700 133.400 101.000 133.700 ;
        RECT 98.900 132.800 99.400 133.100 ;
        RECT 95.800 131.500 96.200 132.500 ;
        RECT 99.000 131.100 99.400 132.800 ;
        RECT 100.600 131.100 101.000 133.400 ;
        RECT 101.400 133.600 103.500 133.900 ;
        RECT 104.000 133.800 105.000 134.200 ;
        RECT 107.000 133.800 108.000 134.200 ;
        RECT 108.300 134.100 109.000 134.500 ;
        RECT 109.400 134.400 109.800 135.200 ;
        RECT 110.200 135.100 110.600 135.200 ;
        RECT 111.000 135.100 111.400 135.200 ;
        RECT 110.200 134.800 111.400 135.100 ;
        RECT 110.200 134.400 110.600 134.800 ;
        RECT 101.400 132.500 101.700 133.600 ;
        RECT 104.000 133.500 104.300 133.800 ;
        RECT 103.900 133.300 104.300 133.500 ;
        RECT 103.500 133.000 104.300 133.300 ;
        RECT 107.700 133.500 108.000 133.800 ;
        RECT 108.500 133.900 109.000 134.100 ;
        RECT 108.500 133.600 110.600 133.900 ;
        RECT 107.700 133.300 108.100 133.500 ;
        RECT 107.700 133.000 108.500 133.300 ;
        RECT 101.400 131.500 101.800 132.500 ;
        RECT 103.500 131.500 103.900 133.000 ;
        RECT 108.100 131.500 108.500 133.000 ;
        RECT 110.300 132.500 110.600 133.600 ;
        RECT 110.200 131.500 110.600 132.500 ;
        RECT 111.000 132.400 111.400 133.200 ;
        RECT 111.800 131.100 112.200 139.900 ;
        RECT 114.500 139.200 114.900 139.900 ;
        RECT 114.500 138.800 115.400 139.200 ;
        RECT 114.500 136.400 114.900 138.800 ;
        RECT 116.600 137.500 117.000 139.500 ;
        RECT 114.100 136.100 114.900 136.400 ;
        RECT 113.400 134.800 113.800 135.600 ;
        RECT 114.100 134.200 114.400 136.100 ;
        RECT 116.700 135.800 117.000 137.500 ;
        RECT 115.100 135.500 117.000 135.800 ;
        RECT 117.400 137.500 117.800 139.500 ;
        RECT 119.500 139.200 119.900 139.900 ;
        RECT 124.100 139.200 124.500 139.900 ;
        RECT 119.500 138.800 120.200 139.200 ;
        RECT 123.800 138.800 124.500 139.200 ;
        RECT 117.400 135.800 117.700 137.500 ;
        RECT 119.500 136.400 119.900 138.800 ;
        RECT 124.100 136.400 124.500 138.800 ;
        RECT 126.200 137.500 126.600 139.500 ;
        RECT 119.500 136.100 120.300 136.400 ;
        RECT 117.400 135.500 119.300 135.800 ;
        RECT 115.100 134.500 115.400 135.500 ;
        RECT 113.400 133.800 114.400 134.200 ;
        RECT 114.700 134.100 115.400 134.500 ;
        RECT 115.800 134.400 116.200 135.200 ;
        RECT 116.600 135.100 117.000 135.200 ;
        RECT 117.400 135.100 117.800 135.200 ;
        RECT 116.600 134.800 117.800 135.100 ;
        RECT 116.600 134.400 117.000 134.800 ;
        RECT 117.400 134.400 117.800 134.800 ;
        RECT 118.200 134.400 118.600 135.200 ;
        RECT 119.000 134.500 119.300 135.500 ;
        RECT 114.100 133.500 114.400 133.800 ;
        RECT 114.900 133.900 115.400 134.100 ;
        RECT 119.000 134.100 119.700 134.500 ;
        RECT 120.000 134.200 120.300 136.100 ;
        RECT 123.700 136.100 124.500 136.400 ;
        RECT 120.600 134.800 121.000 135.600 ;
        RECT 123.000 134.800 123.400 135.600 ;
        RECT 123.700 134.200 124.000 136.100 ;
        RECT 126.300 135.800 126.600 137.500 ;
        RECT 124.700 135.500 126.600 135.800 ;
        RECT 127.000 137.500 127.400 139.500 ;
        RECT 129.100 139.200 129.500 139.900 ;
        RECT 129.100 138.800 129.800 139.200 ;
        RECT 127.000 135.800 127.300 137.500 ;
        RECT 129.100 136.400 129.500 138.800 ;
        RECT 129.100 136.100 129.900 136.400 ;
        RECT 127.000 135.500 128.900 135.800 ;
        RECT 124.700 134.500 125.000 135.500 ;
        RECT 119.000 133.900 119.500 134.100 ;
        RECT 114.900 133.600 117.000 133.900 ;
        RECT 114.100 133.300 114.500 133.500 ;
        RECT 114.100 133.000 114.900 133.300 ;
        RECT 114.500 131.500 114.900 133.000 ;
        RECT 116.700 132.500 117.000 133.600 ;
        RECT 116.600 131.500 117.000 132.500 ;
        RECT 117.400 133.600 119.500 133.900 ;
        RECT 120.000 133.800 121.000 134.200 ;
        RECT 123.000 133.800 124.000 134.200 ;
        RECT 124.300 134.100 125.000 134.500 ;
        RECT 125.400 134.400 125.800 135.200 ;
        RECT 126.200 134.400 126.600 135.200 ;
        RECT 127.000 134.400 127.400 135.200 ;
        RECT 127.800 134.400 128.200 135.200 ;
        RECT 128.600 134.500 128.900 135.500 ;
        RECT 117.400 132.500 117.700 133.600 ;
        RECT 120.000 133.500 120.300 133.800 ;
        RECT 119.900 133.300 120.300 133.500 ;
        RECT 119.500 133.000 120.300 133.300 ;
        RECT 123.700 133.500 124.000 133.800 ;
        RECT 124.500 133.900 125.000 134.100 ;
        RECT 128.600 134.100 129.300 134.500 ;
        RECT 129.600 134.200 129.900 136.100 ;
        RECT 131.800 135.900 132.200 139.900 ;
        RECT 132.600 136.200 133.000 139.900 ;
        RECT 134.200 136.200 134.600 139.900 ;
        RECT 132.600 135.900 134.600 136.200 ;
        RECT 136.300 136.200 136.700 139.900 ;
        RECT 137.000 136.800 137.400 137.200 ;
        RECT 137.100 136.200 137.400 136.800 ;
        RECT 138.500 136.200 138.900 139.900 ;
        RECT 136.300 135.900 136.800 136.200 ;
        RECT 137.100 135.900 137.800 136.200 ;
        RECT 130.200 135.100 130.600 135.600 ;
        RECT 131.900 135.200 132.200 135.900 ;
        RECT 133.800 135.200 134.200 135.400 ;
        RECT 131.000 135.100 131.400 135.200 ;
        RECT 130.200 134.800 131.400 135.100 ;
        RECT 131.800 134.900 133.000 135.200 ;
        RECT 133.800 135.100 134.600 135.200 ;
        RECT 133.800 134.900 135.300 135.100 ;
        RECT 131.800 134.800 132.200 134.900 ;
        RECT 128.600 133.900 129.100 134.100 ;
        RECT 124.500 133.600 126.600 133.900 ;
        RECT 123.700 133.300 124.100 133.500 ;
        RECT 123.700 133.000 124.500 133.300 ;
        RECT 117.400 131.500 117.800 132.500 ;
        RECT 119.500 131.500 119.900 133.000 ;
        RECT 124.100 131.500 124.500 133.000 ;
        RECT 126.300 132.500 126.600 133.600 ;
        RECT 126.200 131.500 126.600 132.500 ;
        RECT 127.000 133.600 129.100 133.900 ;
        RECT 129.600 133.800 130.600 134.200 ;
        RECT 127.000 132.500 127.300 133.600 ;
        RECT 129.600 133.500 129.900 133.800 ;
        RECT 129.500 133.300 129.900 133.500 ;
        RECT 129.100 133.000 129.900 133.300 ;
        RECT 127.000 131.500 127.400 132.500 ;
        RECT 129.100 131.500 129.500 133.000 ;
        RECT 131.800 132.800 132.200 133.200 ;
        RECT 132.700 133.100 133.000 134.900 ;
        RECT 134.200 134.800 135.300 134.900 ;
        RECT 133.400 133.800 133.800 134.600 ;
        RECT 135.000 134.200 135.300 134.800 ;
        RECT 135.800 134.400 136.200 135.200 ;
        RECT 136.500 134.200 136.800 135.900 ;
        RECT 137.400 135.800 137.800 135.900 ;
        RECT 138.200 135.900 138.900 136.200 ;
        RECT 138.200 135.200 138.500 135.900 ;
        RECT 140.600 135.600 141.000 139.900 ;
        RECT 141.400 135.800 141.800 136.600 ;
        RECT 139.000 135.400 141.000 135.600 ;
        RECT 138.900 135.300 141.000 135.400 ;
        RECT 137.400 135.100 137.800 135.200 ;
        RECT 138.200 135.100 138.600 135.200 ;
        RECT 137.400 134.800 138.600 135.100 ;
        RECT 138.900 135.000 139.300 135.300 ;
        RECT 135.000 134.100 135.400 134.200 ;
        RECT 135.000 133.800 135.800 134.100 ;
        RECT 136.500 133.800 137.800 134.200 ;
        RECT 135.400 133.600 135.800 133.800 ;
        RECT 135.100 133.100 136.900 133.300 ;
        RECT 137.400 133.100 137.700 133.800 ;
        RECT 138.200 133.100 138.500 134.800 ;
        RECT 138.900 133.500 139.200 135.000 ;
        RECT 139.600 134.200 140.000 134.600 ;
        RECT 139.700 133.800 140.200 134.200 ;
        RECT 138.900 133.200 140.100 133.500 ;
        RECT 131.900 132.400 132.300 132.800 ;
        RECT 132.600 131.100 133.000 133.100 ;
        RECT 135.000 133.000 137.000 133.100 ;
        RECT 135.000 131.100 135.400 133.000 ;
        RECT 136.600 131.100 137.000 133.000 ;
        RECT 137.400 131.100 137.800 133.100 ;
        RECT 138.200 131.100 138.600 133.100 ;
        RECT 139.800 132.100 140.100 133.200 ;
        RECT 140.600 132.400 141.000 133.200 ;
        RECT 142.200 133.100 142.600 139.900 ;
        RECT 143.000 133.400 143.400 134.200 ;
        RECT 143.800 133.400 144.200 134.200 ;
        RECT 141.700 132.800 142.600 133.100 ;
        RECT 144.600 133.100 145.000 139.900 ;
        RECT 146.600 136.800 147.000 137.200 ;
        RECT 145.400 135.800 145.800 136.600 ;
        RECT 146.600 136.200 146.900 136.800 ;
        RECT 147.300 136.200 147.700 139.900 ;
        RECT 150.200 137.100 150.600 137.200 ;
        RECT 151.800 137.100 152.200 139.900 ;
        RECT 150.200 136.800 152.200 137.100 ;
        RECT 146.200 135.900 146.900 136.200 ;
        RECT 147.200 135.900 147.700 136.200 ;
        RECT 146.200 135.800 146.600 135.900 ;
        RECT 145.400 134.800 145.800 135.200 ;
        RECT 145.400 134.100 145.700 134.800 ;
        RECT 147.200 134.200 147.500 135.900 ;
        RECT 147.800 134.400 148.200 135.200 ;
        RECT 146.200 134.100 147.500 134.200 ;
        RECT 148.600 134.100 149.000 134.200 ;
        RECT 151.800 134.100 152.200 136.800 ;
        RECT 153.900 136.200 154.300 139.900 ;
        RECT 154.600 136.800 155.000 137.200 ;
        RECT 154.700 136.200 155.000 136.800 ;
        RECT 153.900 135.900 154.400 136.200 ;
        RECT 154.700 135.900 155.400 136.200 ;
        RECT 153.400 134.400 153.800 135.200 ;
        RECT 154.100 134.200 154.400 135.900 ;
        RECT 155.000 135.800 155.400 135.900 ;
        RECT 152.600 134.100 153.000 134.200 ;
        RECT 145.400 133.800 147.500 134.100 ;
        RECT 148.200 133.800 150.500 134.100 ;
        RECT 146.300 133.100 146.600 133.800 ;
        RECT 148.200 133.600 148.600 133.800 ;
        RECT 147.100 133.100 148.900 133.300 ;
        RECT 150.200 133.200 150.500 133.800 ;
        RECT 151.800 133.800 153.400 134.100 ;
        RECT 154.100 133.800 155.400 134.200 ;
        RECT 150.200 133.100 150.600 133.200 ;
        RECT 151.000 133.100 151.400 133.200 ;
        RECT 144.600 132.800 145.500 133.100 ;
        RECT 141.700 132.200 142.100 132.800 ;
        RECT 145.100 132.200 145.500 132.800 ;
        RECT 139.800 131.100 140.200 132.100 ;
        RECT 141.700 131.800 142.600 132.200 ;
        RECT 144.600 131.800 145.500 132.200 ;
        RECT 141.700 131.100 142.100 131.800 ;
        RECT 145.100 131.100 145.500 131.800 ;
        RECT 146.200 131.100 146.600 133.100 ;
        RECT 147.000 133.000 149.000 133.100 ;
        RECT 147.000 131.100 147.400 133.000 ;
        RECT 148.600 131.100 149.000 133.000 ;
        RECT 150.200 132.800 151.400 133.100 ;
        RECT 151.000 132.400 151.400 132.800 ;
        RECT 151.800 131.100 152.200 133.800 ;
        RECT 153.000 133.600 153.400 133.800 ;
        RECT 152.700 133.100 154.500 133.300 ;
        RECT 155.000 133.100 155.300 133.800 ;
        RECT 155.800 133.400 156.200 134.200 ;
        RECT 152.600 133.000 154.600 133.100 ;
        RECT 152.600 131.100 153.000 133.000 ;
        RECT 154.200 131.100 154.600 133.000 ;
        RECT 155.000 131.100 155.400 133.100 ;
        RECT 156.600 131.100 157.000 139.900 ;
        RECT 157.400 136.200 157.800 139.900 ;
        RECT 159.000 136.200 159.400 139.900 ;
        RECT 157.400 135.900 159.400 136.200 ;
        RECT 159.800 135.900 160.200 139.900 ;
        RECT 161.900 136.200 162.300 139.900 ;
        RECT 162.600 136.800 163.000 137.200 ;
        RECT 162.700 136.200 163.000 136.800 ;
        RECT 164.200 136.800 164.600 137.200 ;
        RECT 164.200 136.200 164.500 136.800 ;
        RECT 164.900 136.200 165.300 139.900 ;
        RECT 161.900 135.900 162.400 136.200 ;
        RECT 162.700 136.100 163.400 136.200 ;
        RECT 163.800 136.100 164.500 136.200 ;
        RECT 162.700 135.900 164.500 136.100 ;
        RECT 164.800 135.900 165.300 136.200 ;
        RECT 167.000 135.900 167.400 139.900 ;
        RECT 167.800 136.200 168.200 139.900 ;
        RECT 169.400 136.200 169.800 139.900 ;
        RECT 167.800 135.900 169.800 136.200 ;
        RECT 157.800 135.200 158.200 135.400 ;
        RECT 159.800 135.200 160.100 135.900 ;
        RECT 157.400 134.900 158.200 135.200 ;
        RECT 159.000 134.900 160.200 135.200 ;
        RECT 157.400 134.800 157.800 134.900 ;
        RECT 158.200 133.800 158.600 134.600 ;
        RECT 159.000 133.100 159.300 134.900 ;
        RECT 159.800 134.800 160.200 134.900 ;
        RECT 161.400 134.400 161.800 135.200 ;
        RECT 162.100 134.200 162.400 135.900 ;
        RECT 163.000 135.800 164.200 135.900 ;
        RECT 164.800 134.200 165.100 135.900 ;
        RECT 167.100 135.200 167.400 135.900 ;
        RECT 170.200 135.700 170.600 139.900 ;
        RECT 172.400 138.200 172.800 139.900 ;
        RECT 171.800 137.900 172.800 138.200 ;
        RECT 174.600 137.900 175.000 139.900 ;
        RECT 176.700 137.900 177.300 139.900 ;
        RECT 171.800 137.500 172.200 137.900 ;
        RECT 174.600 137.600 174.900 137.900 ;
        RECT 173.500 137.300 175.300 137.600 ;
        RECT 176.600 137.500 177.000 137.900 ;
        RECT 173.500 137.200 173.900 137.300 ;
        RECT 174.900 137.200 175.300 137.300 ;
        RECT 171.800 136.500 172.200 136.600 ;
        RECT 174.100 136.500 174.500 136.600 ;
        RECT 171.800 136.200 174.500 136.500 ;
        RECT 174.800 136.500 175.900 136.800 ;
        RECT 174.800 135.900 175.100 136.500 ;
        RECT 175.500 136.400 175.900 136.500 ;
        RECT 176.700 136.600 177.400 137.000 ;
        RECT 176.700 136.100 177.000 136.600 ;
        RECT 172.700 135.700 175.100 135.900 ;
        RECT 170.200 135.600 175.100 135.700 ;
        RECT 175.800 135.800 177.000 136.100 ;
        RECT 170.200 135.500 173.100 135.600 ;
        RECT 170.200 135.400 173.000 135.500 ;
        RECT 169.000 135.200 169.400 135.400 ;
        RECT 175.800 135.200 176.100 135.800 ;
        RECT 179.000 135.600 179.400 139.900 ;
        RECT 177.300 135.300 179.400 135.600 ;
        RECT 177.300 135.200 177.700 135.300 ;
        RECT 165.400 134.400 165.800 135.200 ;
        RECT 167.000 134.900 168.200 135.200 ;
        RECT 169.000 134.900 169.800 135.200 ;
        RECT 173.400 135.100 173.800 135.200 ;
        RECT 167.000 134.800 167.400 134.900 ;
        RECT 160.600 134.100 161.000 134.200 ;
        RECT 160.600 133.800 161.400 134.100 ;
        RECT 162.100 133.800 163.400 134.200 ;
        RECT 163.800 133.800 165.100 134.200 ;
        RECT 166.200 134.100 166.600 134.200 ;
        RECT 165.800 133.800 166.600 134.100 ;
        RECT 167.000 134.100 167.400 134.200 ;
        RECT 167.900 134.100 168.200 134.900 ;
        RECT 169.400 134.800 169.800 134.900 ;
        RECT 171.300 134.800 173.800 135.100 ;
        RECT 175.800 134.800 176.200 135.200 ;
        RECT 178.100 134.900 178.500 135.000 ;
        RECT 171.300 134.700 171.700 134.800 ;
        RECT 172.600 134.700 173.000 134.800 ;
        RECT 167.000 133.800 168.200 134.100 ;
        RECT 168.600 133.800 169.000 134.600 ;
        RECT 172.100 134.200 172.500 134.300 ;
        RECT 175.800 134.200 176.100 134.800 ;
        RECT 176.600 134.600 178.500 134.900 ;
        RECT 176.600 134.500 177.000 134.600 ;
        RECT 170.600 133.900 176.100 134.200 ;
        RECT 170.600 133.800 171.400 133.900 ;
        RECT 161.000 133.600 161.400 133.800 ;
        RECT 159.000 131.100 159.400 133.100 ;
        RECT 159.800 132.800 160.200 133.200 ;
        RECT 160.700 133.100 162.500 133.300 ;
        RECT 163.000 133.100 163.300 133.800 ;
        RECT 163.900 133.100 164.200 133.800 ;
        RECT 165.800 133.600 166.200 133.800 ;
        RECT 164.700 133.100 166.500 133.300 ;
        RECT 160.600 133.000 162.600 133.100 ;
        RECT 159.700 132.400 160.100 132.800 ;
        RECT 160.600 131.100 161.000 133.000 ;
        RECT 162.200 131.100 162.600 133.000 ;
        RECT 163.000 131.100 163.400 133.100 ;
        RECT 163.800 131.100 164.200 133.100 ;
        RECT 164.600 133.000 166.600 133.100 ;
        RECT 164.600 131.100 165.000 133.000 ;
        RECT 166.200 131.100 166.600 133.000 ;
        RECT 167.000 132.800 167.400 133.200 ;
        RECT 167.900 133.100 168.200 133.800 ;
        RECT 167.100 132.400 167.500 132.800 ;
        RECT 167.800 131.100 168.200 133.100 ;
        RECT 170.200 131.100 170.600 133.500 ;
        RECT 172.700 132.800 173.000 133.900 ;
        RECT 175.500 133.800 175.900 133.900 ;
        RECT 179.000 133.600 179.400 135.300 ;
        RECT 177.500 133.300 179.400 133.600 ;
        RECT 177.500 133.200 177.900 133.300 ;
        RECT 171.800 132.100 172.200 132.500 ;
        RECT 172.600 132.400 173.000 132.800 ;
        RECT 173.500 132.700 173.900 132.800 ;
        RECT 173.500 132.400 174.900 132.700 ;
        RECT 174.600 132.100 174.900 132.400 ;
        RECT 176.600 132.100 177.000 132.500 ;
        RECT 179.000 132.100 179.400 133.300 ;
        RECT 179.800 135.600 180.200 139.900 ;
        RECT 181.900 137.900 182.500 139.900 ;
        RECT 184.200 137.900 184.600 139.900 ;
        RECT 186.400 138.200 186.800 139.900 ;
        RECT 186.400 137.900 187.400 138.200 ;
        RECT 182.200 137.500 182.600 137.900 ;
        RECT 184.300 137.600 184.600 137.900 ;
        RECT 183.900 137.300 185.700 137.600 ;
        RECT 187.000 137.500 187.400 137.900 ;
        RECT 183.900 137.200 184.300 137.300 ;
        RECT 185.300 137.200 185.700 137.300 ;
        RECT 181.800 136.600 182.500 137.000 ;
        RECT 182.200 136.100 182.500 136.600 ;
        RECT 183.300 136.500 184.400 136.800 ;
        RECT 183.300 136.400 183.700 136.500 ;
        RECT 182.200 135.800 183.400 136.100 ;
        RECT 179.800 135.300 181.900 135.600 ;
        RECT 179.800 133.600 180.200 135.300 ;
        RECT 181.500 135.200 181.900 135.300 ;
        RECT 183.100 135.200 183.400 135.800 ;
        RECT 184.100 135.900 184.400 136.500 ;
        RECT 184.700 136.500 185.100 136.600 ;
        RECT 187.000 136.500 187.400 136.600 ;
        RECT 184.700 136.200 187.400 136.500 ;
        RECT 184.100 135.700 186.500 135.900 ;
        RECT 188.600 135.700 189.000 139.900 ;
        RECT 189.400 136.200 189.800 139.900 ;
        RECT 191.800 136.200 192.200 139.900 ;
        RECT 189.400 135.900 190.500 136.200 ;
        RECT 191.800 135.900 192.900 136.200 ;
        RECT 184.100 135.600 189.000 135.700 ;
        RECT 186.100 135.500 189.000 135.600 ;
        RECT 186.200 135.400 189.000 135.500 ;
        RECT 190.200 135.600 190.500 135.900 ;
        RECT 192.600 135.600 192.900 135.900 ;
        RECT 190.200 135.200 190.800 135.600 ;
        RECT 192.600 135.200 193.200 135.600 ;
        RECT 180.700 134.900 181.100 135.000 ;
        RECT 180.700 134.600 182.600 134.900 ;
        RECT 183.000 134.800 183.400 135.200 ;
        RECT 183.800 135.100 184.200 135.200 ;
        RECT 185.400 135.100 185.800 135.200 ;
        RECT 183.800 134.800 187.900 135.100 ;
        RECT 182.200 134.500 182.600 134.600 ;
        RECT 183.100 134.200 183.400 134.800 ;
        RECT 187.500 134.700 187.900 134.800 ;
        RECT 186.700 134.200 187.100 134.300 ;
        RECT 183.100 133.900 188.600 134.200 ;
        RECT 183.300 133.800 183.700 133.900 ;
        RECT 179.800 133.300 181.700 133.600 ;
        RECT 179.800 132.100 180.200 133.300 ;
        RECT 181.300 133.200 181.700 133.300 ;
        RECT 186.200 132.800 186.500 133.900 ;
        RECT 187.800 133.800 188.600 133.900 ;
        RECT 190.200 133.700 190.500 135.200 ;
        RECT 191.800 134.400 192.200 135.200 ;
        RECT 192.600 133.700 192.900 135.200 ;
        RECT 185.300 132.700 185.700 132.800 ;
        RECT 182.200 132.100 182.600 132.500 ;
        RECT 184.300 132.400 185.700 132.700 ;
        RECT 186.200 132.400 186.600 132.800 ;
        RECT 184.300 132.100 184.600 132.400 ;
        RECT 187.000 132.100 187.400 132.500 ;
        RECT 171.800 131.800 172.800 132.100 ;
        RECT 172.400 131.100 172.800 131.800 ;
        RECT 174.600 131.100 175.000 132.100 ;
        RECT 176.600 131.800 177.300 132.100 ;
        RECT 176.700 131.100 177.300 131.800 ;
        RECT 179.000 131.800 180.200 132.100 ;
        RECT 179.000 131.100 179.400 131.800 ;
        RECT 179.800 131.100 180.200 131.800 ;
        RECT 181.900 131.800 182.600 132.100 ;
        RECT 181.900 131.100 182.500 131.800 ;
        RECT 184.200 131.100 184.600 132.100 ;
        RECT 186.400 131.800 187.400 132.100 ;
        RECT 186.400 131.100 186.800 131.800 ;
        RECT 188.600 131.100 189.000 133.500 ;
        RECT 189.400 133.400 190.500 133.700 ;
        RECT 191.800 133.400 192.900 133.700 ;
        RECT 189.400 131.100 189.800 133.400 ;
        RECT 191.800 131.100 192.200 133.400 ;
        RECT 0.600 127.700 1.000 129.900 ;
        RECT 2.700 129.200 3.300 129.900 ;
        RECT 2.700 128.900 3.400 129.200 ;
        RECT 5.000 128.900 5.400 129.900 ;
        RECT 7.200 129.200 7.600 129.900 ;
        RECT 7.200 128.900 8.200 129.200 ;
        RECT 3.000 128.500 3.400 128.900 ;
        RECT 5.100 128.600 5.400 128.900 ;
        RECT 5.100 128.300 6.500 128.600 ;
        RECT 6.100 128.200 6.500 128.300 ;
        RECT 7.000 128.200 7.400 128.600 ;
        RECT 7.800 128.500 8.200 128.900 ;
        RECT 2.100 127.700 2.500 127.800 ;
        RECT 0.600 127.400 2.500 127.700 ;
        RECT 0.600 125.700 1.000 127.400 ;
        RECT 4.100 127.100 4.500 127.200 ;
        RECT 7.000 127.100 7.300 128.200 ;
        RECT 9.400 127.500 9.800 129.900 ;
        RECT 10.200 127.700 10.600 129.900 ;
        RECT 12.300 129.200 12.900 129.900 ;
        RECT 12.300 128.900 13.000 129.200 ;
        RECT 14.600 128.900 15.000 129.900 ;
        RECT 16.800 129.200 17.200 129.900 ;
        RECT 16.800 128.900 17.800 129.200 ;
        RECT 12.600 128.500 13.000 128.900 ;
        RECT 14.700 128.600 15.000 128.900 ;
        RECT 14.700 128.300 16.100 128.600 ;
        RECT 15.700 128.200 16.100 128.300 ;
        RECT 16.600 128.200 17.000 128.600 ;
        RECT 17.400 128.500 17.800 128.900 ;
        RECT 11.700 127.700 12.100 127.800 ;
        RECT 10.200 127.400 12.100 127.700 ;
        RECT 8.600 127.100 9.400 127.200 ;
        RECT 3.900 126.800 9.400 127.100 ;
        RECT 3.000 126.400 3.400 126.500 ;
        RECT 1.500 126.100 3.400 126.400 ;
        RECT 1.500 126.000 1.900 126.100 ;
        RECT 2.300 125.700 2.700 125.800 ;
        RECT 0.600 125.400 2.700 125.700 ;
        RECT 0.600 121.100 1.000 125.400 ;
        RECT 3.900 125.200 4.200 126.800 ;
        RECT 7.500 126.700 7.900 126.800 ;
        RECT 8.300 126.200 8.700 126.300 ;
        RECT 6.200 125.900 8.700 126.200 ;
        RECT 6.200 125.800 6.600 125.900 ;
        RECT 10.200 125.700 10.600 127.400 ;
        RECT 11.000 126.800 11.400 127.400 ;
        RECT 13.700 127.100 14.600 127.200 ;
        RECT 16.600 127.100 16.900 128.200 ;
        RECT 19.000 127.500 19.400 129.900 ;
        RECT 19.800 127.500 20.200 129.900 ;
        RECT 22.000 129.200 22.400 129.900 ;
        RECT 21.400 128.900 22.400 129.200 ;
        RECT 24.200 128.900 24.600 129.900 ;
        RECT 26.300 129.200 26.900 129.900 ;
        RECT 26.200 128.900 26.900 129.200 ;
        RECT 21.400 128.500 21.800 128.900 ;
        RECT 24.200 128.600 24.500 128.900 ;
        RECT 22.200 128.200 22.600 128.600 ;
        RECT 23.100 128.300 24.500 128.600 ;
        RECT 26.200 128.500 26.600 128.900 ;
        RECT 23.100 128.200 23.500 128.300 ;
        RECT 18.200 127.100 19.000 127.200 ;
        RECT 13.500 126.800 19.000 127.100 ;
        RECT 20.200 127.100 21.000 127.200 ;
        RECT 22.300 127.100 22.600 128.200 ;
        RECT 27.100 127.700 27.500 127.800 ;
        RECT 28.600 127.700 29.000 129.900 ;
        RECT 27.100 127.400 29.000 127.700 ;
        RECT 25.100 127.100 25.500 127.200 ;
        RECT 20.200 126.800 25.700 127.100 ;
        RECT 12.600 126.400 13.000 126.500 ;
        RECT 11.100 126.100 13.000 126.400 ;
        RECT 11.100 126.000 11.500 126.100 ;
        RECT 11.900 125.700 12.300 125.800 ;
        RECT 7.000 125.500 9.800 125.600 ;
        RECT 6.900 125.400 9.800 125.500 ;
        RECT 3.000 124.900 4.200 125.200 ;
        RECT 4.900 125.300 9.800 125.400 ;
        RECT 4.900 125.100 7.300 125.300 ;
        RECT 3.000 124.400 3.300 124.900 ;
        RECT 2.600 124.000 3.300 124.400 ;
        RECT 4.100 124.500 4.500 124.600 ;
        RECT 4.900 124.500 5.200 125.100 ;
        RECT 4.100 124.200 5.200 124.500 ;
        RECT 5.500 124.500 8.200 124.800 ;
        RECT 5.500 124.400 5.900 124.500 ;
        RECT 7.800 124.400 8.200 124.500 ;
        RECT 4.700 123.700 5.100 123.800 ;
        RECT 6.100 123.700 6.500 123.800 ;
        RECT 3.000 123.100 3.400 123.500 ;
        RECT 4.700 123.400 6.500 123.700 ;
        RECT 5.100 123.100 5.400 123.400 ;
        RECT 7.800 123.100 8.200 123.500 ;
        RECT 2.700 121.100 3.300 123.100 ;
        RECT 5.000 121.100 5.400 123.100 ;
        RECT 7.200 122.800 8.200 123.100 ;
        RECT 7.200 121.100 7.600 122.800 ;
        RECT 9.400 121.100 9.800 125.300 ;
        RECT 10.200 125.400 12.300 125.700 ;
        RECT 10.200 121.100 10.600 125.400 ;
        RECT 13.500 125.200 13.800 126.800 ;
        RECT 17.100 126.700 17.500 126.800 ;
        RECT 21.700 126.700 22.100 126.800 ;
        RECT 16.600 126.200 17.000 126.300 ;
        RECT 17.900 126.200 18.300 126.300 ;
        RECT 15.800 125.900 18.300 126.200 ;
        RECT 20.900 126.200 21.300 126.300 ;
        RECT 25.400 126.200 25.700 126.800 ;
        RECT 26.200 126.400 26.600 126.500 ;
        RECT 20.900 126.100 23.400 126.200 ;
        RECT 23.800 126.100 24.200 126.200 ;
        RECT 20.900 125.900 24.200 126.100 ;
        RECT 15.800 125.800 16.200 125.900 ;
        RECT 23.000 125.800 24.200 125.900 ;
        RECT 25.400 125.800 25.800 126.200 ;
        RECT 26.200 126.100 28.100 126.400 ;
        RECT 27.700 126.000 28.100 126.100 ;
        RECT 16.600 125.500 19.400 125.600 ;
        RECT 16.500 125.400 19.400 125.500 ;
        RECT 12.600 124.900 13.800 125.200 ;
        RECT 14.500 125.300 19.400 125.400 ;
        RECT 14.500 125.100 16.900 125.300 ;
        RECT 12.600 124.400 12.900 124.900 ;
        RECT 12.200 124.000 12.900 124.400 ;
        RECT 13.700 124.500 14.100 124.600 ;
        RECT 14.500 124.500 14.800 125.100 ;
        RECT 13.700 124.200 14.800 124.500 ;
        RECT 15.100 124.500 17.800 124.800 ;
        RECT 15.100 124.400 15.500 124.500 ;
        RECT 17.400 124.400 17.800 124.500 ;
        RECT 14.300 123.700 14.700 123.800 ;
        RECT 15.700 123.700 16.100 123.800 ;
        RECT 12.600 123.100 13.000 123.500 ;
        RECT 14.300 123.400 16.100 123.700 ;
        RECT 14.700 123.100 15.000 123.400 ;
        RECT 17.400 123.100 17.800 123.500 ;
        RECT 12.300 121.100 12.900 123.100 ;
        RECT 14.600 121.100 15.000 123.100 ;
        RECT 16.800 122.800 17.800 123.100 ;
        RECT 16.800 121.100 17.200 122.800 ;
        RECT 19.000 121.100 19.400 125.300 ;
        RECT 19.800 125.500 22.600 125.600 ;
        RECT 19.800 125.400 22.700 125.500 ;
        RECT 19.800 125.300 24.700 125.400 ;
        RECT 19.800 121.100 20.200 125.300 ;
        RECT 22.300 125.100 24.700 125.300 ;
        RECT 21.400 124.500 24.100 124.800 ;
        RECT 21.400 124.400 21.800 124.500 ;
        RECT 23.700 124.400 24.100 124.500 ;
        RECT 24.400 124.500 24.700 125.100 ;
        RECT 25.400 125.200 25.700 125.800 ;
        RECT 26.900 125.700 27.300 125.800 ;
        RECT 28.600 125.700 29.000 127.400 ;
        RECT 29.400 126.800 29.800 127.600 ;
        RECT 29.400 126.200 29.700 126.800 ;
        RECT 29.400 125.800 29.800 126.200 ;
        RECT 26.900 125.400 29.000 125.700 ;
        RECT 25.400 124.900 26.600 125.200 ;
        RECT 25.100 124.500 25.500 124.600 ;
        RECT 24.400 124.200 25.500 124.500 ;
        RECT 26.300 124.400 26.600 124.900 ;
        RECT 26.300 124.000 27.000 124.400 ;
        RECT 23.100 123.700 23.500 123.800 ;
        RECT 24.500 123.700 24.900 123.800 ;
        RECT 21.400 123.100 21.800 123.500 ;
        RECT 23.100 123.400 24.900 123.700 ;
        RECT 24.200 123.100 24.500 123.400 ;
        RECT 26.200 123.100 26.600 123.500 ;
        RECT 21.400 122.800 22.400 123.100 ;
        RECT 22.000 121.100 22.400 122.800 ;
        RECT 24.200 121.100 24.600 123.100 ;
        RECT 26.300 121.100 26.900 123.100 ;
        RECT 28.600 121.100 29.000 125.400 ;
        RECT 30.200 121.100 30.600 129.900 ;
        RECT 32.300 128.200 32.700 129.900 ;
        RECT 31.800 127.900 32.700 128.200 ;
        RECT 31.000 126.800 31.400 127.600 ;
        RECT 31.800 126.100 32.200 127.900 ;
        RECT 33.400 127.800 33.800 128.600 ;
        RECT 32.600 126.100 33.000 126.200 ;
        RECT 31.800 125.800 33.000 126.100 ;
        RECT 31.800 121.100 32.200 125.800 ;
        RECT 32.600 125.100 33.000 125.200 ;
        RECT 33.400 125.100 33.800 125.200 ;
        RECT 32.600 124.800 33.800 125.100 ;
        RECT 34.200 125.100 34.600 129.900 ;
        RECT 35.000 127.900 35.400 129.900 ;
        RECT 35.800 128.000 36.200 129.900 ;
        RECT 37.400 128.000 37.800 129.900 ;
        RECT 39.000 128.900 39.400 129.900 ;
        RECT 35.800 127.900 37.800 128.000 ;
        RECT 35.100 127.200 35.400 127.900 ;
        RECT 35.900 127.700 37.700 127.900 ;
        RECT 38.200 127.800 38.600 128.600 ;
        RECT 37.000 127.200 37.400 127.400 ;
        RECT 39.100 127.200 39.400 128.900 ;
        RECT 35.000 126.800 36.300 127.200 ;
        RECT 37.000 126.900 37.800 127.200 ;
        RECT 37.400 126.800 37.800 126.900 ;
        RECT 39.000 126.800 39.400 127.200 ;
        RECT 41.200 127.100 41.600 129.900 ;
        RECT 43.800 127.800 44.200 128.600 ;
        RECT 35.000 125.100 35.400 125.200 ;
        RECT 36.000 125.100 36.300 126.800 ;
        RECT 36.600 126.100 37.000 126.600 ;
        RECT 37.400 126.100 37.800 126.200 ;
        RECT 36.600 125.800 37.800 126.100 ;
        RECT 39.100 125.100 39.400 126.800 ;
        RECT 40.700 126.900 41.600 127.100 ;
        RECT 40.700 126.800 41.500 126.900 ;
        RECT 39.800 125.400 40.200 126.200 ;
        RECT 40.700 125.200 41.000 126.800 ;
        RECT 41.800 125.800 42.600 126.200 ;
        RECT 34.200 124.800 35.700 125.100 ;
        RECT 36.000 124.800 36.500 125.100 ;
        RECT 32.600 124.400 33.000 124.800 ;
        RECT 34.200 121.100 34.600 124.800 ;
        RECT 35.400 124.200 35.700 124.800 ;
        RECT 35.400 123.800 35.800 124.200 ;
        RECT 36.100 122.200 36.500 124.800 ;
        RECT 39.000 124.700 39.900 125.100 ;
        RECT 40.600 124.800 41.000 125.200 ;
        RECT 43.000 124.800 43.400 125.600 ;
        RECT 44.600 125.100 45.000 129.900 ;
        RECT 45.400 129.100 45.800 129.200 ;
        RECT 47.000 129.100 47.400 129.900 ;
        RECT 45.400 128.800 47.400 129.100 ;
        RECT 47.000 127.900 47.400 128.800 ;
        RECT 47.800 128.000 48.200 129.900 ;
        RECT 49.400 128.000 49.800 129.900 ;
        RECT 47.800 127.900 49.800 128.000 ;
        RECT 51.000 128.800 51.400 129.900 ;
        RECT 47.100 127.200 47.400 127.900 ;
        RECT 47.900 127.700 49.700 127.900 ;
        RECT 49.000 127.200 49.400 127.400 ;
        RECT 51.000 127.200 51.300 128.800 ;
        RECT 51.800 127.800 52.200 128.600 ;
        RECT 52.600 127.800 53.000 128.600 ;
        RECT 47.000 126.800 48.300 127.200 ;
        RECT 49.000 126.900 49.800 127.200 ;
        RECT 49.400 126.800 49.800 126.900 ;
        RECT 51.000 126.800 51.400 127.200 ;
        RECT 47.000 125.100 47.400 125.200 ;
        RECT 48.000 125.100 48.300 126.800 ;
        RECT 48.600 125.800 49.000 126.600 ;
        RECT 50.200 125.400 50.600 126.200 ;
        RECT 51.000 125.100 51.300 126.800 ;
        RECT 53.400 125.100 53.800 129.900 ;
        RECT 56.000 127.100 56.400 129.900 ;
        RECT 58.200 128.900 58.600 129.900 ;
        RECT 57.400 127.800 57.800 128.600 ;
        RECT 58.300 127.200 58.600 128.900 ;
        RECT 60.100 128.200 60.500 129.900 ;
        RECT 62.500 128.200 62.900 129.900 ;
        RECT 65.200 129.200 65.600 129.900 ;
        RECT 65.200 128.800 65.800 129.200 ;
        RECT 68.600 128.900 69.000 129.900 ;
        RECT 71.800 129.200 72.200 129.900 ;
        RECT 59.000 128.100 59.400 128.200 ;
        RECT 60.100 128.100 61.000 128.200 ;
        RECT 59.000 127.800 61.000 128.100 ;
        RECT 62.500 127.900 63.400 128.200 ;
        RECT 56.000 126.900 56.900 127.100 ;
        RECT 56.100 126.800 56.900 126.900 ;
        RECT 58.200 126.800 58.600 127.200 ;
        RECT 55.000 125.800 55.800 126.200 ;
        RECT 54.200 125.100 54.600 125.600 ;
        RECT 44.600 124.800 47.700 125.100 ;
        RECT 48.000 124.800 48.500 125.100 ;
        RECT 39.500 124.200 39.900 124.700 ;
        RECT 39.500 123.800 40.200 124.200 ;
        RECT 36.100 121.800 37.000 122.200 ;
        RECT 36.100 121.100 36.500 121.800 ;
        RECT 39.500 121.100 39.900 123.800 ;
        RECT 40.700 123.500 41.000 124.800 ;
        RECT 41.400 123.800 41.800 124.600 ;
        RECT 40.700 123.200 42.500 123.500 ;
        RECT 40.700 123.100 41.000 123.200 ;
        RECT 40.600 121.100 41.000 123.100 ;
        RECT 42.200 121.100 42.600 123.200 ;
        RECT 44.600 121.100 45.000 124.800 ;
        RECT 47.400 124.200 47.700 124.800 ;
        RECT 47.400 123.800 47.800 124.200 ;
        RECT 48.100 121.100 48.500 124.800 ;
        RECT 50.500 124.700 51.400 125.100 ;
        RECT 53.400 124.800 54.600 125.100 ;
        RECT 56.600 125.200 56.900 126.800 ;
        RECT 56.600 124.800 57.000 125.200 ;
        RECT 58.300 125.100 58.600 126.800 ;
        RECT 59.000 126.100 59.400 126.200 ;
        RECT 59.000 125.800 60.100 126.100 ;
        RECT 59.000 125.400 59.400 125.800 ;
        RECT 59.800 125.200 60.100 125.800 ;
        RECT 50.500 122.200 50.900 124.700 ;
        RECT 50.200 121.800 50.900 122.200 ;
        RECT 50.500 121.100 50.900 121.800 ;
        RECT 53.400 121.100 53.800 124.800 ;
        RECT 55.800 123.800 56.200 124.600 ;
        RECT 56.600 123.500 56.900 124.800 ;
        RECT 58.200 124.700 59.100 125.100 ;
        RECT 58.700 124.200 59.100 124.700 ;
        RECT 59.800 124.400 60.200 125.200 ;
        RECT 58.200 123.800 59.100 124.200 ;
        RECT 55.100 123.200 56.900 123.500 ;
        RECT 55.100 123.100 55.400 123.200 ;
        RECT 55.000 121.100 55.400 123.100 ;
        RECT 56.600 123.100 56.900 123.200 ;
        RECT 56.600 121.100 57.000 123.100 ;
        RECT 58.700 121.100 59.100 123.800 ;
        RECT 60.600 121.100 61.000 127.800 ;
        RECT 61.400 126.800 61.800 127.600 ;
        RECT 61.400 125.100 61.800 125.200 ;
        RECT 62.200 125.100 62.600 125.200 ;
        RECT 61.400 124.800 62.600 125.100 ;
        RECT 62.200 124.400 62.600 124.800 ;
        RECT 63.000 121.100 63.400 127.900 ;
        RECT 63.800 126.800 64.200 127.600 ;
        RECT 65.200 127.100 65.600 128.800 ;
        RECT 68.600 127.200 68.900 128.900 ;
        RECT 71.800 128.800 72.300 129.200 ;
        RECT 73.400 128.900 73.800 129.900 ;
        RECT 77.400 128.900 77.800 129.900 ;
        RECT 73.400 128.800 74.000 128.900 ;
        RECT 69.400 128.100 69.800 128.600 ;
        RECT 72.000 128.500 74.000 128.800 ;
        RECT 71.000 128.100 71.900 128.200 ;
        RECT 72.600 128.100 73.000 128.200 ;
        RECT 69.400 127.800 73.000 128.100 ;
        RECT 64.700 126.900 65.600 127.100 ;
        RECT 67.800 127.100 68.200 127.200 ;
        RECT 68.600 127.100 69.000 127.200 ;
        RECT 64.700 126.800 65.500 126.900 ;
        RECT 67.800 126.800 69.000 127.100 ;
        RECT 71.800 126.800 72.600 127.200 ;
        RECT 64.700 125.200 65.000 126.800 ;
        RECT 65.800 125.800 66.600 126.200 ;
        RECT 64.600 124.800 65.000 125.200 ;
        RECT 67.000 124.800 67.400 125.600 ;
        RECT 67.800 125.400 68.200 126.200 ;
        RECT 68.600 125.100 68.900 126.800 ;
        RECT 72.600 125.800 73.400 126.200 ;
        RECT 73.700 125.200 74.000 128.500 ;
        RECT 76.600 127.800 77.000 128.600 ;
        RECT 77.500 127.200 77.800 128.900 ;
        RECT 79.000 128.000 79.400 129.900 ;
        RECT 80.600 128.000 81.000 129.900 ;
        RECT 79.000 127.900 81.000 128.000 ;
        RECT 81.400 127.900 81.800 129.900 ;
        RECT 82.500 129.200 82.900 129.900 ;
        RECT 82.200 128.800 82.900 129.200 ;
        RECT 82.500 128.200 82.900 128.800 ;
        RECT 82.500 127.900 83.400 128.200 ;
        RECT 79.100 127.700 80.900 127.900 ;
        RECT 79.400 127.200 79.800 127.400 ;
        RECT 81.400 127.200 81.700 127.900 ;
        RECT 77.400 126.800 77.800 127.200 ;
        RECT 78.200 127.100 78.600 127.200 ;
        RECT 79.000 127.100 79.800 127.200 ;
        RECT 78.200 126.900 79.800 127.100 ;
        RECT 78.200 126.800 79.400 126.900 ;
        RECT 80.500 126.800 81.800 127.200 ;
        RECT 64.700 123.500 65.000 124.800 ;
        RECT 68.100 124.700 69.000 125.100 ;
        RECT 73.700 124.900 75.400 125.200 ;
        RECT 77.500 125.100 77.800 126.800 ;
        RECT 78.200 126.100 78.600 126.200 ;
        RECT 79.800 126.100 80.200 126.600 ;
        RECT 78.200 125.800 80.200 126.100 ;
        RECT 78.200 125.400 78.600 125.800 ;
        RECT 80.500 125.200 80.800 126.800 ;
        RECT 75.000 124.800 75.400 124.900 ;
        RECT 65.400 123.800 65.800 124.600 ;
        RECT 64.700 123.200 66.500 123.500 ;
        RECT 64.700 123.100 65.000 123.200 ;
        RECT 64.600 121.100 65.000 123.100 ;
        RECT 66.200 123.100 66.500 123.200 ;
        RECT 66.200 121.100 66.600 123.100 ;
        RECT 68.100 121.100 68.500 124.700 ;
        RECT 70.300 124.400 72.100 124.700 ;
        RECT 70.300 124.100 70.600 124.400 ;
        RECT 70.200 121.100 70.600 124.100 ;
        RECT 71.800 124.100 72.100 124.400 ;
        RECT 72.700 124.500 74.500 124.600 ;
        RECT 75.000 124.500 75.300 124.800 ;
        RECT 77.400 124.700 78.300 125.100 ;
        RECT 79.800 124.800 80.800 125.200 ;
        RECT 81.400 125.100 81.800 125.200 ;
        RECT 82.200 125.100 82.600 125.200 ;
        RECT 81.100 124.800 82.600 125.100 ;
        RECT 72.700 124.300 74.600 124.500 ;
        RECT 72.700 124.100 73.000 124.300 ;
        RECT 71.800 121.400 72.200 124.100 ;
        RECT 72.600 121.700 73.000 124.100 ;
        RECT 73.400 121.400 73.800 124.000 ;
        RECT 74.200 121.500 74.600 124.300 ;
        RECT 75.000 121.700 75.400 124.500 ;
        RECT 71.800 121.100 73.800 121.400 ;
        RECT 74.300 121.400 74.600 121.500 ;
        RECT 75.800 121.500 76.200 124.500 ;
        RECT 77.900 124.200 78.300 124.700 ;
        RECT 77.400 123.800 78.300 124.200 ;
        RECT 75.800 121.400 76.100 121.500 ;
        RECT 74.300 121.100 76.100 121.400 ;
        RECT 77.900 121.100 78.300 123.800 ;
        RECT 80.300 121.100 80.700 124.800 ;
        RECT 81.100 124.200 81.400 124.800 ;
        RECT 82.200 124.400 82.600 124.800 ;
        RECT 81.000 123.800 81.400 124.200 ;
        RECT 83.000 121.100 83.400 127.900 ;
        RECT 83.800 127.100 84.200 127.600 ;
        RECT 84.600 127.100 85.000 127.600 ;
        RECT 83.800 126.800 85.000 127.100 ;
        RECT 85.400 127.100 85.800 129.900 ;
        RECT 87.800 128.800 88.200 129.900 ;
        RECT 87.000 127.800 87.400 128.600 ;
        RECT 87.000 127.100 87.300 127.800 ;
        RECT 87.900 127.200 88.200 128.800 ;
        RECT 85.400 126.800 87.300 127.100 ;
        RECT 87.800 126.800 88.200 127.200 ;
        RECT 84.600 126.100 85.000 126.200 ;
        RECT 85.400 126.100 85.800 126.800 ;
        RECT 84.600 125.800 85.800 126.100 ;
        RECT 85.400 121.100 85.800 125.800 ;
        RECT 87.900 125.100 88.200 126.800 ;
        RECT 88.600 126.100 89.000 126.200 ;
        RECT 89.400 126.100 89.800 129.900 ;
        RECT 90.200 128.100 90.600 128.600 ;
        RECT 91.000 128.100 91.400 129.900 ;
        RECT 93.100 129.200 93.700 129.900 ;
        RECT 93.100 128.900 93.800 129.200 ;
        RECT 95.400 128.900 95.800 129.900 ;
        RECT 97.600 129.200 98.000 129.900 ;
        RECT 97.600 128.900 98.600 129.200 ;
        RECT 93.400 128.500 93.800 128.900 ;
        RECT 95.500 128.600 95.800 128.900 ;
        RECT 95.500 128.300 96.900 128.600 ;
        RECT 96.500 128.200 96.900 128.300 ;
        RECT 97.400 128.200 97.800 128.600 ;
        RECT 98.200 128.500 98.600 128.900 ;
        RECT 90.200 127.800 91.400 128.100 ;
        RECT 88.600 125.800 89.800 126.100 ;
        RECT 88.600 125.400 89.000 125.800 ;
        RECT 87.800 124.700 88.700 125.100 ;
        RECT 88.300 121.100 88.700 124.700 ;
        RECT 89.400 121.100 89.800 125.800 ;
        RECT 91.000 127.700 91.400 127.800 ;
        RECT 92.500 127.700 92.900 127.800 ;
        RECT 91.000 127.400 92.900 127.700 ;
        RECT 91.000 125.700 91.400 127.400 ;
        RECT 94.500 127.100 94.900 127.200 ;
        RECT 97.400 127.100 97.700 128.200 ;
        RECT 99.800 127.500 100.200 129.900 ;
        RECT 103.000 127.600 103.400 129.900 ;
        RECT 104.600 127.600 105.000 129.900 ;
        RECT 106.200 127.600 106.600 129.900 ;
        RECT 107.800 127.600 108.200 129.900 ;
        RECT 110.200 128.200 110.600 129.900 ;
        RECT 102.200 127.200 103.400 127.600 ;
        RECT 103.900 127.200 105.000 127.600 ;
        RECT 105.500 127.200 106.600 127.600 ;
        RECT 107.300 127.200 108.200 127.600 ;
        RECT 110.100 127.900 110.600 128.200 ;
        RECT 110.100 127.200 110.400 127.900 ;
        RECT 111.800 127.600 112.200 129.900 ;
        RECT 110.900 127.300 112.200 127.600 ;
        RECT 112.600 128.500 113.000 129.500 ;
        RECT 112.600 127.400 112.900 128.500 ;
        RECT 114.700 128.000 115.100 129.500 ;
        RECT 114.700 127.700 115.500 128.000 ;
        RECT 117.400 127.800 117.800 128.600 ;
        RECT 115.100 127.500 115.500 127.700 ;
        RECT 99.000 127.100 99.800 127.200 ;
        RECT 94.300 126.800 99.800 127.100 ;
        RECT 93.400 126.400 93.800 126.500 ;
        RECT 91.900 126.100 93.800 126.400 ;
        RECT 91.900 126.000 92.300 126.100 ;
        RECT 92.700 125.700 93.100 125.800 ;
        RECT 91.000 125.400 93.100 125.700 ;
        RECT 91.000 121.100 91.400 125.400 ;
        RECT 94.300 125.200 94.600 126.800 ;
        RECT 97.900 126.700 98.300 126.800 ;
        RECT 98.700 126.200 99.100 126.300 ;
        RECT 96.600 125.900 99.100 126.200 ;
        RECT 96.600 125.800 97.000 125.900 ;
        RECT 102.200 125.800 102.600 127.200 ;
        RECT 103.900 126.900 104.300 127.200 ;
        RECT 105.500 126.900 105.900 127.200 ;
        RECT 107.300 126.900 107.700 127.200 ;
        RECT 103.000 126.500 104.300 126.900 ;
        RECT 104.700 126.500 105.900 126.900 ;
        RECT 106.400 126.500 107.700 126.900 ;
        RECT 103.900 125.800 104.300 126.500 ;
        RECT 105.500 125.800 105.900 126.500 ;
        RECT 107.300 125.800 107.700 126.500 ;
        RECT 110.100 126.800 110.600 127.200 ;
        RECT 97.400 125.500 100.200 125.600 ;
        RECT 97.300 125.400 100.200 125.500 ;
        RECT 102.200 125.400 103.400 125.800 ;
        RECT 103.900 125.400 105.000 125.800 ;
        RECT 105.500 125.400 106.600 125.800 ;
        RECT 107.300 125.400 108.200 125.800 ;
        RECT 93.400 124.900 94.600 125.200 ;
        RECT 95.300 125.300 100.200 125.400 ;
        RECT 95.300 125.100 97.700 125.300 ;
        RECT 93.400 124.400 93.700 124.900 ;
        RECT 93.000 124.000 93.700 124.400 ;
        RECT 94.500 124.500 94.900 124.600 ;
        RECT 95.300 124.500 95.600 125.100 ;
        RECT 94.500 124.200 95.600 124.500 ;
        RECT 95.900 124.500 98.600 124.800 ;
        RECT 95.900 124.400 96.300 124.500 ;
        RECT 98.200 124.400 98.600 124.500 ;
        RECT 95.100 123.700 95.500 123.800 ;
        RECT 96.500 123.700 96.900 123.800 ;
        RECT 93.400 123.100 93.800 123.500 ;
        RECT 95.100 123.400 96.900 123.700 ;
        RECT 95.500 123.100 95.800 123.400 ;
        RECT 98.200 123.100 98.600 123.500 ;
        RECT 93.100 121.100 93.700 123.100 ;
        RECT 95.400 121.100 95.800 123.100 ;
        RECT 97.600 122.800 98.600 123.100 ;
        RECT 97.600 121.100 98.000 122.800 ;
        RECT 99.800 121.100 100.200 125.300 ;
        RECT 103.000 121.100 103.400 125.400 ;
        RECT 104.600 121.100 105.000 125.400 ;
        RECT 106.200 121.100 106.600 125.400 ;
        RECT 107.800 121.100 108.200 125.400 ;
        RECT 110.100 125.100 110.400 126.800 ;
        RECT 110.900 126.500 111.200 127.300 ;
        RECT 112.600 127.100 114.700 127.400 ;
        RECT 114.200 126.900 114.700 127.100 ;
        RECT 115.200 127.200 115.500 127.500 ;
        RECT 110.700 126.100 111.200 126.500 ;
        RECT 110.900 125.100 111.200 126.100 ;
        RECT 111.700 126.200 112.100 126.600 ;
        RECT 111.700 125.800 112.200 126.200 ;
        RECT 112.600 125.800 113.000 126.600 ;
        RECT 113.400 125.800 113.800 126.600 ;
        RECT 114.200 126.500 114.900 126.900 ;
        RECT 115.200 126.800 116.200 127.200 ;
        RECT 114.200 125.500 114.500 126.500 ;
        RECT 112.600 125.200 114.500 125.500 ;
        RECT 110.100 124.600 110.600 125.100 ;
        RECT 110.900 124.800 112.200 125.100 ;
        RECT 110.200 121.100 110.600 124.600 ;
        RECT 111.800 121.100 112.200 124.800 ;
        RECT 112.600 123.500 112.900 125.200 ;
        RECT 115.200 124.900 115.500 126.800 ;
        RECT 115.800 125.400 116.200 126.200 ;
        RECT 114.700 124.600 115.500 124.900 ;
        RECT 112.600 121.500 113.000 123.500 ;
        RECT 114.700 122.200 115.100 124.600 ;
        RECT 114.700 121.800 115.400 122.200 ;
        RECT 114.700 121.100 115.100 121.800 ;
        RECT 118.200 121.100 118.600 129.900 ;
        RECT 119.800 128.200 120.200 129.900 ;
        RECT 119.700 127.800 120.200 128.200 ;
        RECT 119.700 127.200 120.000 127.800 ;
        RECT 121.400 127.600 121.800 129.900 ;
        RECT 120.500 127.300 121.800 127.600 ;
        RECT 123.000 127.600 123.400 129.900 ;
        RECT 124.600 127.600 125.000 129.900 ;
        RECT 126.200 127.600 126.600 129.900 ;
        RECT 127.800 127.600 128.200 129.900 ;
        RECT 129.400 127.600 129.800 129.900 ;
        RECT 131.000 128.200 131.400 129.900 ;
        RECT 131.000 127.900 131.500 128.200 ;
        RECT 119.700 126.800 120.200 127.200 ;
        RECT 119.700 125.100 120.000 126.800 ;
        RECT 120.500 126.500 120.800 127.300 ;
        RECT 123.000 127.200 123.900 127.600 ;
        RECT 124.600 127.200 125.700 127.600 ;
        RECT 126.200 127.200 127.300 127.600 ;
        RECT 127.800 127.200 129.000 127.600 ;
        RECT 129.400 127.300 130.700 127.600 ;
        RECT 123.500 126.900 123.900 127.200 ;
        RECT 125.300 126.900 125.700 127.200 ;
        RECT 126.900 126.900 127.300 127.200 ;
        RECT 120.300 126.100 120.800 126.500 ;
        RECT 120.500 125.100 120.800 126.100 ;
        RECT 121.300 126.200 121.700 126.600 ;
        RECT 123.500 126.500 124.800 126.900 ;
        RECT 125.300 126.500 126.500 126.900 ;
        RECT 126.900 126.500 128.200 126.900 ;
        RECT 121.300 126.100 121.800 126.200 ;
        RECT 122.200 126.100 122.600 126.200 ;
        RECT 121.300 125.800 122.600 126.100 ;
        RECT 123.500 125.800 123.900 126.500 ;
        RECT 125.300 125.800 125.700 126.500 ;
        RECT 126.900 125.800 127.300 126.500 ;
        RECT 128.600 125.800 129.000 127.200 ;
        RECT 129.500 126.200 129.900 126.600 ;
        RECT 129.400 125.800 129.900 126.200 ;
        RECT 130.400 126.500 130.700 127.300 ;
        RECT 131.200 127.200 131.500 127.900 ;
        RECT 132.600 127.600 133.000 129.900 ;
        RECT 134.200 128.200 134.600 129.900 ;
        RECT 134.200 127.900 134.700 128.200 ;
        RECT 132.600 127.300 133.900 127.600 ;
        RECT 131.000 126.800 131.500 127.200 ;
        RECT 130.400 126.100 130.900 126.500 ;
        RECT 123.000 125.400 123.900 125.800 ;
        RECT 124.600 125.400 125.700 125.800 ;
        RECT 126.200 125.400 127.300 125.800 ;
        RECT 127.800 125.400 129.000 125.800 ;
        RECT 119.700 124.600 120.200 125.100 ;
        RECT 120.500 124.800 121.800 125.100 ;
        RECT 119.800 121.100 120.200 124.600 ;
        RECT 121.400 121.100 121.800 124.800 ;
        RECT 123.000 121.100 123.400 125.400 ;
        RECT 124.600 121.100 125.000 125.400 ;
        RECT 126.200 121.100 126.600 125.400 ;
        RECT 127.800 121.100 128.200 125.400 ;
        RECT 130.400 125.100 130.700 126.100 ;
        RECT 131.200 125.100 131.500 126.800 ;
        RECT 132.700 126.200 133.100 126.600 ;
        RECT 132.600 125.800 133.100 126.200 ;
        RECT 133.600 126.500 133.900 127.300 ;
        RECT 134.400 127.200 134.700 127.900 ;
        RECT 134.200 126.800 134.700 127.200 ;
        RECT 135.000 127.100 135.400 127.200 ;
        RECT 135.800 127.100 136.200 129.900 ;
        RECT 137.400 128.000 137.800 129.900 ;
        RECT 139.000 128.000 139.400 129.900 ;
        RECT 137.400 127.900 139.400 128.000 ;
        RECT 139.800 128.100 140.200 129.900 ;
        RECT 140.700 128.200 141.100 128.600 ;
        RECT 140.600 128.100 141.000 128.200 ;
        RECT 137.500 127.700 139.300 127.900 ;
        RECT 139.800 127.800 141.000 128.100 ;
        RECT 141.400 127.900 141.800 129.900 ;
        RECT 145.100 128.200 145.500 129.900 ;
        RECT 147.000 128.800 147.400 129.900 ;
        RECT 135.000 126.800 136.200 127.100 ;
        RECT 136.600 126.800 137.000 127.600 ;
        RECT 137.800 127.200 138.200 127.400 ;
        RECT 139.800 127.200 140.100 127.800 ;
        RECT 137.400 126.900 138.200 127.200 ;
        RECT 137.400 126.800 137.800 126.900 ;
        RECT 138.900 126.800 140.200 127.200 ;
        RECT 133.600 126.100 134.100 126.500 ;
        RECT 133.600 125.100 133.900 126.100 ;
        RECT 134.400 125.100 134.700 126.800 ;
        RECT 129.400 124.800 130.700 125.100 ;
        RECT 129.400 121.100 129.800 124.800 ;
        RECT 131.000 124.600 131.500 125.100 ;
        RECT 132.600 124.800 133.900 125.100 ;
        RECT 131.000 121.100 131.400 124.600 ;
        RECT 132.600 121.100 133.000 124.800 ;
        RECT 134.200 124.600 134.700 125.100 ;
        RECT 134.200 121.100 134.600 124.600 ;
        RECT 135.800 121.100 136.200 126.800 ;
        RECT 138.200 125.800 138.600 126.600 ;
        RECT 138.900 125.100 139.200 126.800 ;
        RECT 141.500 126.200 141.800 127.900 ;
        RECT 144.600 128.100 145.500 128.200 ;
        RECT 146.200 128.100 146.600 128.600 ;
        RECT 144.600 127.800 146.600 128.100 ;
        RECT 142.200 126.400 142.600 127.200 ;
        RECT 143.800 126.800 144.200 127.600 ;
        RECT 140.600 126.100 141.000 126.200 ;
        RECT 141.400 126.100 141.800 126.200 ;
        RECT 143.000 126.100 143.400 126.200 ;
        RECT 140.600 125.800 141.800 126.100 ;
        RECT 142.600 125.800 143.400 126.100 ;
        RECT 144.600 126.100 145.000 127.800 ;
        RECT 147.100 127.200 147.400 128.800 ;
        RECT 147.000 126.800 147.400 127.200 ;
        RECT 145.400 126.100 145.800 126.200 ;
        RECT 144.600 125.800 145.800 126.100 ;
        RECT 139.800 125.100 140.200 125.200 ;
        RECT 140.700 125.100 141.000 125.800 ;
        RECT 142.600 125.600 143.000 125.800 ;
        RECT 138.700 124.800 139.200 125.100 ;
        RECT 139.500 124.800 140.200 125.100 ;
        RECT 138.700 121.100 139.100 124.800 ;
        RECT 139.500 124.200 139.800 124.800 ;
        RECT 139.400 123.800 139.800 124.200 ;
        RECT 140.600 121.100 141.000 125.100 ;
        RECT 141.400 124.800 143.400 125.100 ;
        RECT 141.400 121.100 141.800 124.800 ;
        RECT 143.000 121.100 143.400 124.800 ;
        RECT 144.600 121.100 145.000 125.800 ;
        RECT 145.400 124.400 145.800 125.200 ;
        RECT 147.100 125.100 147.400 126.800 ;
        RECT 151.000 128.900 151.400 129.900 ;
        RECT 151.000 127.200 151.300 128.900 ;
        RECT 151.800 127.800 152.200 128.600 ;
        RECT 154.200 127.900 154.600 129.900 ;
        RECT 154.900 128.200 155.300 128.600 ;
        RECT 151.000 127.100 151.400 127.200 ;
        RECT 153.400 127.100 153.800 127.200 ;
        RECT 151.000 126.800 153.800 127.100 ;
        RECT 147.800 125.400 148.200 126.200 ;
        RECT 150.200 125.400 150.600 126.200 ;
        RECT 151.000 125.100 151.300 126.800 ;
        RECT 153.400 126.400 153.800 126.800 ;
        RECT 152.600 126.100 153.000 126.200 ;
        RECT 154.200 126.100 154.500 127.900 ;
        RECT 155.000 127.800 155.400 128.200 ;
        RECT 155.000 126.800 155.400 127.200 ;
        RECT 156.400 127.100 156.800 129.900 ;
        RECT 159.300 128.200 159.700 129.900 ;
        RECT 162.200 128.900 162.600 129.900 ;
        RECT 155.900 126.900 156.800 127.100 ;
        RECT 159.000 127.800 160.200 128.200 ;
        RECT 159.000 127.200 159.300 127.800 ;
        RECT 155.900 126.800 156.700 126.900 ;
        RECT 159.000 126.800 159.400 127.200 ;
        RECT 155.000 126.200 155.300 126.800 ;
        RECT 155.000 126.100 155.400 126.200 ;
        RECT 152.600 125.800 153.400 126.100 ;
        RECT 154.200 125.800 155.400 126.100 ;
        RECT 153.000 125.600 153.400 125.800 ;
        RECT 155.000 125.100 155.300 125.800 ;
        RECT 155.900 125.200 156.200 126.800 ;
        RECT 157.000 125.800 157.800 126.200 ;
        RECT 147.000 124.700 147.900 125.100 ;
        RECT 147.500 121.100 147.900 124.700 ;
        RECT 150.500 124.700 151.400 125.100 ;
        RECT 152.600 124.800 154.600 125.100 ;
        RECT 150.500 122.200 150.900 124.700 ;
        RECT 150.200 121.800 150.900 122.200 ;
        RECT 150.500 121.100 150.900 121.800 ;
        RECT 152.600 121.100 153.000 124.800 ;
        RECT 154.200 121.100 154.600 124.800 ;
        RECT 155.000 121.100 155.400 125.100 ;
        RECT 155.800 124.800 156.200 125.200 ;
        RECT 158.200 124.800 158.600 125.600 ;
        RECT 155.900 123.500 156.200 124.800 ;
        RECT 156.600 123.800 157.000 124.600 ;
        RECT 157.400 124.100 157.800 124.200 ;
        RECT 159.000 124.100 159.400 125.200 ;
        RECT 157.400 123.800 159.400 124.100 ;
        RECT 155.900 123.200 157.700 123.500 ;
        RECT 155.900 123.100 156.200 123.200 ;
        RECT 155.800 121.100 156.200 123.100 ;
        RECT 157.400 123.100 157.700 123.200 ;
        RECT 157.400 121.100 157.800 123.100 ;
        RECT 159.800 121.100 160.200 127.800 ;
        RECT 160.600 126.800 161.000 127.600 ;
        RECT 162.200 127.200 162.500 128.900 ;
        RECT 163.000 128.100 163.400 128.600 ;
        RECT 163.800 128.100 164.200 129.900 ;
        RECT 163.000 127.800 164.200 128.100 ;
        RECT 164.600 128.000 165.000 129.900 ;
        RECT 166.200 128.000 166.600 129.900 ;
        RECT 164.600 127.900 166.600 128.000 ;
        RECT 167.000 127.900 167.400 129.900 ;
        RECT 169.200 129.200 170.000 129.900 ;
        RECT 168.600 128.800 170.000 129.200 ;
        RECT 169.200 128.100 170.000 128.800 ;
        RECT 163.900 127.200 164.200 127.800 ;
        RECT 164.700 127.700 166.500 127.900 ;
        RECT 167.000 127.600 168.200 127.900 ;
        RECT 167.800 127.500 168.200 127.600 ;
        RECT 168.500 127.400 168.900 127.800 ;
        RECT 165.800 127.200 166.200 127.400 ;
        RECT 168.500 127.200 168.800 127.400 ;
        RECT 162.200 126.800 162.600 127.200 ;
        RECT 163.000 126.800 163.400 127.200 ;
        RECT 163.800 126.800 165.100 127.200 ;
        RECT 165.800 126.900 166.600 127.200 ;
        RECT 166.200 126.800 166.600 126.900 ;
        RECT 167.000 126.800 167.800 127.200 ;
        RECT 168.400 126.800 168.800 127.200 ;
        RECT 161.400 125.400 161.800 126.200 ;
        RECT 162.200 126.100 162.500 126.800 ;
        RECT 163.000 126.100 163.300 126.800 ;
        RECT 162.200 125.800 163.300 126.100 ;
        RECT 162.200 125.100 162.500 125.800 ;
        RECT 163.800 125.100 164.200 125.200 ;
        RECT 164.800 125.100 165.100 126.800 ;
        RECT 165.400 125.800 165.800 126.600 ;
        RECT 169.200 126.400 169.500 128.100 ;
        RECT 171.800 127.900 172.200 129.900 ;
        RECT 169.800 127.700 170.600 127.800 ;
        RECT 169.800 127.400 170.800 127.700 ;
        RECT 171.100 127.600 172.200 127.900 ;
        RECT 172.600 127.700 173.000 129.900 ;
        RECT 174.700 129.200 175.300 129.900 ;
        RECT 174.700 128.900 175.400 129.200 ;
        RECT 177.000 128.900 177.400 129.900 ;
        RECT 179.200 129.200 179.600 129.900 ;
        RECT 179.200 128.900 180.200 129.200 ;
        RECT 175.000 128.500 175.400 128.900 ;
        RECT 177.100 128.600 177.400 128.900 ;
        RECT 177.100 128.300 178.500 128.600 ;
        RECT 178.100 128.200 178.500 128.300 ;
        RECT 179.000 128.200 179.400 128.600 ;
        RECT 179.800 128.500 180.200 128.900 ;
        RECT 174.100 127.700 174.500 127.800 ;
        RECT 171.100 127.500 171.500 127.600 ;
        RECT 170.500 127.200 170.800 127.400 ;
        RECT 172.600 127.400 174.500 127.700 ;
        RECT 169.800 126.700 170.200 127.100 ;
        RECT 170.500 126.900 172.200 127.200 ;
        RECT 171.400 126.800 172.200 126.900 ;
        RECT 169.000 126.200 169.500 126.400 ;
        RECT 168.600 126.100 169.500 126.200 ;
        RECT 169.900 126.400 170.200 126.700 ;
        RECT 169.900 126.100 171.200 126.400 ;
        RECT 168.600 125.800 169.300 126.100 ;
        RECT 170.800 126.000 171.200 126.100 ;
        RECT 169.000 125.100 169.300 125.800 ;
        RECT 169.700 125.700 170.100 125.800 ;
        RECT 172.600 125.700 173.000 127.400 ;
        RECT 176.100 127.100 176.500 127.200 ;
        RECT 179.000 127.100 179.300 128.200 ;
        RECT 181.400 127.500 181.800 129.900 ;
        RECT 184.100 128.200 184.500 129.500 ;
        RECT 186.200 128.500 186.600 129.500 ;
        RECT 184.100 128.000 185.000 128.200 ;
        RECT 183.700 127.800 185.000 128.000 ;
        RECT 183.700 127.700 184.500 127.800 ;
        RECT 183.700 127.500 184.100 127.700 ;
        RECT 183.700 127.200 184.000 127.500 ;
        RECT 186.300 127.400 186.600 128.500 ;
        RECT 187.000 127.800 187.400 128.600 ;
        RECT 180.600 127.100 181.400 127.200 ;
        RECT 175.900 126.800 181.400 127.100 ;
        RECT 183.000 126.800 184.000 127.200 ;
        RECT 184.500 127.100 186.600 127.400 ;
        RECT 184.500 126.900 185.000 127.100 ;
        RECT 175.000 126.400 175.400 126.500 ;
        RECT 173.500 126.100 175.400 126.400 ;
        RECT 175.900 126.200 176.200 126.800 ;
        RECT 179.500 126.700 179.900 126.800 ;
        RECT 180.300 126.200 180.700 126.300 ;
        RECT 173.500 126.000 173.900 126.100 ;
        RECT 175.800 125.800 176.200 126.200 ;
        RECT 178.200 125.900 180.700 126.200 ;
        RECT 178.200 125.800 178.600 125.900 ;
        RECT 174.300 125.700 174.700 125.800 ;
        RECT 169.700 125.400 171.400 125.700 ;
        RECT 171.100 125.100 171.400 125.400 ;
        RECT 172.600 125.400 174.700 125.700 ;
        RECT 161.700 124.700 162.600 125.100 ;
        RECT 163.800 124.800 164.500 125.100 ;
        RECT 164.800 124.800 165.300 125.100 ;
        RECT 161.700 121.100 162.100 124.700 ;
        RECT 164.200 124.200 164.500 124.800 ;
        RECT 164.200 123.800 164.600 124.200 ;
        RECT 164.900 121.100 165.300 124.800 ;
        RECT 167.000 124.800 168.200 125.100 ;
        RECT 169.000 124.800 170.000 125.100 ;
        RECT 167.000 121.100 167.400 124.800 ;
        RECT 167.800 124.700 168.200 124.800 ;
        RECT 169.200 121.100 170.000 124.800 ;
        RECT 171.100 124.800 172.200 125.100 ;
        RECT 171.100 124.700 171.500 124.800 ;
        RECT 171.800 121.100 172.200 124.800 ;
        RECT 172.600 121.100 173.000 125.400 ;
        RECT 175.900 125.200 176.200 125.800 ;
        RECT 179.000 125.500 181.800 125.600 ;
        RECT 178.900 125.400 181.800 125.500 ;
        RECT 183.000 125.400 183.400 126.200 ;
        RECT 175.000 124.900 176.200 125.200 ;
        RECT 176.900 125.300 181.800 125.400 ;
        RECT 176.900 125.100 179.300 125.300 ;
        RECT 175.000 124.400 175.300 124.900 ;
        RECT 174.600 124.200 175.300 124.400 ;
        RECT 176.100 124.500 176.500 124.600 ;
        RECT 176.900 124.500 177.200 125.100 ;
        RECT 176.100 124.200 177.200 124.500 ;
        RECT 177.500 124.500 180.200 124.800 ;
        RECT 177.500 124.400 177.900 124.500 ;
        RECT 179.800 124.400 180.200 124.500 ;
        RECT 174.200 124.000 175.300 124.200 ;
        RECT 174.200 123.800 174.900 124.000 ;
        RECT 176.700 123.700 177.100 123.800 ;
        RECT 178.100 123.700 178.500 123.800 ;
        RECT 175.000 123.100 175.400 123.500 ;
        RECT 176.700 123.400 178.500 123.700 ;
        RECT 177.100 123.100 177.400 123.400 ;
        RECT 179.800 123.100 180.200 123.500 ;
        RECT 174.700 121.100 175.300 123.100 ;
        RECT 177.000 121.100 177.400 123.100 ;
        RECT 179.200 122.800 180.200 123.100 ;
        RECT 179.200 121.100 179.600 122.800 ;
        RECT 181.400 121.100 181.800 125.300 ;
        RECT 183.700 124.900 184.000 126.800 ;
        RECT 184.300 126.500 185.000 126.900 ;
        RECT 184.700 125.500 185.000 126.500 ;
        RECT 185.400 125.800 185.800 126.600 ;
        RECT 186.200 125.800 186.600 126.600 ;
        RECT 184.700 125.200 186.600 125.500 ;
        RECT 183.700 124.600 184.500 124.900 ;
        RECT 184.100 121.100 184.500 124.600 ;
        RECT 186.300 123.500 186.600 125.200 ;
        RECT 186.200 121.500 186.600 123.500 ;
        RECT 187.800 121.100 188.200 129.900 ;
        RECT 189.400 128.900 189.800 129.900 ;
        RECT 188.600 127.800 189.000 128.600 ;
        RECT 189.500 127.200 189.800 128.900 ;
        RECT 191.000 127.600 191.400 129.900 ;
        RECT 194.200 128.900 194.600 129.900 ;
        RECT 193.400 127.800 193.800 128.600 ;
        RECT 191.000 127.300 192.100 127.600 ;
        RECT 189.400 126.800 189.800 127.200 ;
        RECT 189.500 126.200 189.800 126.800 ;
        RECT 189.400 125.800 189.800 126.200 ;
        RECT 189.500 125.100 189.800 125.800 ;
        RECT 190.200 125.400 190.600 126.200 ;
        RECT 191.000 125.800 191.400 126.600 ;
        RECT 191.800 125.800 192.100 127.300 ;
        RECT 194.300 127.200 194.600 128.900 ;
        RECT 194.200 126.800 194.600 127.200 ;
        RECT 191.800 125.400 192.400 125.800 ;
        RECT 191.800 125.100 192.100 125.400 ;
        RECT 194.300 125.100 194.600 126.800 ;
        RECT 195.000 125.400 195.400 126.200 ;
        RECT 189.400 124.700 190.300 125.100 ;
        RECT 189.900 121.100 190.300 124.700 ;
        RECT 191.000 124.800 192.100 125.100 ;
        RECT 191.000 121.100 191.400 124.800 ;
        RECT 194.200 124.700 195.100 125.100 ;
        RECT 194.700 122.200 195.100 124.700 ;
        RECT 194.700 121.800 195.400 122.200 ;
        RECT 194.700 121.100 195.100 121.800 ;
        RECT 0.600 115.600 1.000 119.900 ;
        RECT 2.700 117.900 3.300 119.900 ;
        RECT 5.000 117.900 5.400 119.900 ;
        RECT 7.200 118.200 7.600 119.900 ;
        RECT 7.200 117.900 8.200 118.200 ;
        RECT 3.000 117.500 3.400 117.900 ;
        RECT 5.100 117.600 5.400 117.900 ;
        RECT 4.700 117.300 6.500 117.600 ;
        RECT 7.800 117.500 8.200 117.900 ;
        RECT 4.700 117.200 5.100 117.300 ;
        RECT 6.100 117.200 6.500 117.300 ;
        RECT 2.600 116.600 3.300 117.000 ;
        RECT 3.000 116.100 3.300 116.600 ;
        RECT 4.100 116.500 5.200 116.800 ;
        RECT 4.100 116.400 4.500 116.500 ;
        RECT 3.000 115.800 4.200 116.100 ;
        RECT 0.600 115.300 2.700 115.600 ;
        RECT 0.600 113.600 1.000 115.300 ;
        RECT 2.300 115.200 2.700 115.300 ;
        RECT 1.500 114.900 1.900 115.000 ;
        RECT 1.500 114.600 3.400 114.900 ;
        RECT 3.000 114.500 3.400 114.600 ;
        RECT 3.900 114.200 4.200 115.800 ;
        RECT 4.900 115.900 5.200 116.500 ;
        RECT 5.500 116.500 5.900 116.600 ;
        RECT 7.800 116.500 8.200 116.600 ;
        RECT 5.500 116.200 8.200 116.500 ;
        RECT 4.900 115.700 7.300 115.900 ;
        RECT 9.400 115.700 9.800 119.900 ;
        RECT 11.500 116.300 11.900 119.900 ;
        RECT 13.400 117.900 13.800 119.900 ;
        RECT 11.000 115.900 11.900 116.300 ;
        RECT 4.900 115.600 9.800 115.700 ;
        RECT 6.900 115.500 9.800 115.600 ;
        RECT 7.000 115.400 9.800 115.500 ;
        RECT 6.200 115.100 6.600 115.200 ;
        RECT 6.200 114.800 8.700 115.100 ;
        RECT 8.300 114.700 8.700 114.800 ;
        RECT 7.500 114.200 7.900 114.300 ;
        RECT 11.100 114.200 11.400 115.900 ;
        RECT 13.500 115.800 13.800 117.900 ;
        RECT 15.000 115.900 15.400 119.900 ;
        RECT 11.800 114.800 12.200 115.600 ;
        RECT 13.500 115.500 14.700 115.800 ;
        RECT 13.400 114.800 13.800 115.200 ;
        RECT 3.900 113.900 9.400 114.200 ;
        RECT 4.100 113.800 4.500 113.900 ;
        RECT 7.000 113.800 7.400 113.900 ;
        RECT 8.600 113.800 9.400 113.900 ;
        RECT 11.000 113.800 11.400 114.200 ;
        RECT 12.600 113.800 13.000 114.600 ;
        RECT 13.500 114.400 13.800 114.800 ;
        RECT 13.400 114.000 14.000 114.400 ;
        RECT 14.400 113.800 14.700 115.500 ;
        RECT 15.100 115.200 15.400 115.900 ;
        RECT 15.800 115.700 16.200 119.900 ;
        RECT 18.000 118.200 18.400 119.900 ;
        RECT 17.400 117.900 18.400 118.200 ;
        RECT 20.200 117.900 20.600 119.900 ;
        RECT 22.300 117.900 22.900 119.900 ;
        RECT 24.600 119.100 25.000 119.900 ;
        RECT 25.400 119.100 25.800 119.900 ;
        RECT 24.600 118.800 25.800 119.100 ;
        RECT 17.400 117.500 17.800 117.900 ;
        RECT 20.200 117.600 20.500 117.900 ;
        RECT 19.100 117.300 20.900 117.600 ;
        RECT 22.200 117.500 22.600 117.900 ;
        RECT 19.100 117.200 19.500 117.300 ;
        RECT 20.500 117.200 20.900 117.300 ;
        RECT 17.400 116.500 17.800 116.600 ;
        RECT 19.700 116.500 20.100 116.600 ;
        RECT 17.400 116.200 20.100 116.500 ;
        RECT 20.400 116.500 21.500 116.800 ;
        RECT 20.400 115.900 20.700 116.500 ;
        RECT 21.100 116.400 21.500 116.500 ;
        RECT 22.300 116.600 23.000 117.000 ;
        RECT 22.300 116.100 22.600 116.600 ;
        RECT 18.300 115.700 20.700 115.900 ;
        RECT 15.800 115.600 20.700 115.700 ;
        RECT 21.400 115.800 22.600 116.100 ;
        RECT 15.800 115.500 18.700 115.600 ;
        RECT 15.800 115.400 18.600 115.500 ;
        RECT 15.000 114.800 15.400 115.200 ;
        RECT 19.000 115.100 19.400 115.200 ;
        RECT 0.600 113.300 2.500 113.600 ;
        RECT 0.600 111.100 1.000 113.300 ;
        RECT 2.100 113.200 2.500 113.300 ;
        RECT 7.000 112.800 7.300 113.800 ;
        RECT 6.100 112.700 6.500 112.800 ;
        RECT 3.000 112.100 3.400 112.500 ;
        RECT 5.100 112.400 6.500 112.700 ;
        RECT 7.000 112.400 7.400 112.800 ;
        RECT 5.100 112.100 5.400 112.400 ;
        RECT 7.800 112.100 8.200 112.500 ;
        RECT 2.700 111.800 3.400 112.100 ;
        RECT 2.700 111.100 3.300 111.800 ;
        RECT 5.000 111.100 5.400 112.100 ;
        RECT 7.200 111.800 8.200 112.100 ;
        RECT 7.200 111.100 7.600 111.800 ;
        RECT 9.400 111.100 9.800 113.500 ;
        RECT 10.200 112.400 10.600 113.200 ;
        RECT 11.100 112.200 11.400 113.800 ;
        RECT 14.400 113.700 14.800 113.800 ;
        RECT 13.300 113.500 14.800 113.700 ;
        RECT 12.700 113.400 14.800 113.500 ;
        RECT 12.700 113.200 13.600 113.400 ;
        RECT 12.700 113.100 13.000 113.200 ;
        RECT 15.100 113.100 15.400 114.800 ;
        RECT 16.900 114.800 19.400 115.100 ;
        RECT 16.900 114.700 17.300 114.800 ;
        RECT 17.700 114.200 18.100 114.300 ;
        RECT 21.400 114.200 21.700 115.800 ;
        RECT 24.600 115.600 25.000 118.800 ;
        RECT 22.900 115.300 25.000 115.600 ;
        RECT 22.900 115.200 23.300 115.300 ;
        RECT 23.700 114.900 24.100 115.000 ;
        RECT 22.200 114.600 24.100 114.900 ;
        RECT 22.200 114.500 22.600 114.600 ;
        RECT 16.200 113.900 21.700 114.200 ;
        RECT 16.200 113.800 17.000 113.900 ;
        RECT 11.000 111.100 11.400 112.200 ;
        RECT 12.600 111.100 13.000 113.100 ;
        RECT 14.700 112.600 15.400 113.100 ;
        RECT 14.700 112.200 15.100 112.600 ;
        RECT 14.700 111.800 15.400 112.200 ;
        RECT 14.700 111.100 15.100 111.800 ;
        RECT 15.800 111.100 16.200 113.500 ;
        RECT 18.300 113.200 18.600 113.900 ;
        RECT 21.100 113.800 21.500 113.900 ;
        RECT 24.600 113.600 25.000 115.300 ;
        RECT 23.100 113.300 25.000 113.600 ;
        RECT 23.100 113.200 23.500 113.300 ;
        RECT 17.400 112.100 17.800 112.500 ;
        RECT 18.200 112.400 18.600 113.200 ;
        RECT 19.100 112.700 19.500 112.800 ;
        RECT 19.100 112.400 20.500 112.700 ;
        RECT 20.200 112.100 20.500 112.400 ;
        RECT 22.200 112.100 22.600 112.500 ;
        RECT 17.400 111.800 18.400 112.100 ;
        RECT 18.000 111.100 18.400 111.800 ;
        RECT 20.200 111.100 20.600 112.100 ;
        RECT 22.200 111.800 22.900 112.100 ;
        RECT 22.300 111.100 22.900 111.800 ;
        RECT 24.600 111.100 25.000 113.300 ;
        RECT 25.400 115.600 25.800 118.800 ;
        RECT 27.500 117.900 28.100 119.900 ;
        RECT 29.800 117.900 30.200 119.900 ;
        RECT 32.000 118.200 32.400 119.900 ;
        RECT 32.000 117.900 33.000 118.200 ;
        RECT 27.800 117.500 28.200 117.900 ;
        RECT 29.900 117.600 30.200 117.900 ;
        RECT 29.500 117.300 31.300 117.600 ;
        RECT 32.600 117.500 33.000 117.900 ;
        RECT 29.500 117.200 29.900 117.300 ;
        RECT 30.900 117.200 31.300 117.300 ;
        RECT 27.400 116.600 28.100 117.000 ;
        RECT 27.800 116.100 28.100 116.600 ;
        RECT 28.900 116.500 30.000 116.800 ;
        RECT 28.900 116.400 29.300 116.500 ;
        RECT 27.800 115.800 29.000 116.100 ;
        RECT 25.400 115.300 27.500 115.600 ;
        RECT 25.400 113.600 25.800 115.300 ;
        RECT 27.100 115.200 27.500 115.300 ;
        RECT 28.700 115.200 29.000 115.800 ;
        RECT 29.700 115.900 30.000 116.500 ;
        RECT 30.300 116.500 30.700 116.600 ;
        RECT 32.600 116.500 33.000 116.600 ;
        RECT 30.300 116.200 33.000 116.500 ;
        RECT 29.700 115.700 32.100 115.900 ;
        RECT 34.200 115.700 34.600 119.900 ;
        RECT 36.300 116.200 36.700 119.900 ;
        RECT 37.000 116.800 37.400 117.200 ;
        RECT 37.100 116.200 37.400 116.800 ;
        RECT 36.300 115.900 36.800 116.200 ;
        RECT 37.100 115.900 37.800 116.200 ;
        RECT 38.200 115.900 38.600 119.900 ;
        RECT 39.000 116.200 39.400 119.900 ;
        RECT 40.600 116.200 41.000 119.900 ;
        RECT 42.700 117.200 43.100 119.900 ;
        RECT 43.800 117.900 44.200 119.900 ;
        RECT 43.900 117.800 44.200 117.900 ;
        RECT 45.400 117.900 45.800 119.900 ;
        RECT 48.600 117.900 49.000 119.900 ;
        RECT 45.400 117.800 45.700 117.900 ;
        RECT 43.900 117.500 45.700 117.800 ;
        RECT 48.700 117.800 49.000 117.900 ;
        RECT 50.200 117.900 50.600 119.900 ;
        RECT 50.200 117.800 50.500 117.900 ;
        RECT 51.800 117.800 52.200 119.900 ;
        RECT 53.400 117.900 53.800 119.900 ;
        RECT 53.400 117.800 53.700 117.900 ;
        RECT 48.700 117.500 50.500 117.800 ;
        RECT 42.700 116.800 43.400 117.200 ;
        RECT 42.700 116.300 43.100 116.800 ;
        RECT 39.000 115.900 41.000 116.200 ;
        RECT 42.200 115.900 43.100 116.300 ;
        RECT 43.900 116.200 44.200 117.500 ;
        RECT 44.600 116.400 45.000 117.200 ;
        RECT 48.700 116.200 49.000 117.500 ;
        RECT 49.400 116.400 49.800 117.200 ;
        RECT 50.200 117.100 50.500 117.500 ;
        RECT 51.900 117.500 53.700 117.800 ;
        RECT 51.000 117.100 51.400 117.200 ;
        RECT 50.200 116.800 51.400 117.100 ;
        RECT 51.900 116.200 52.200 117.500 ;
        RECT 52.600 116.400 53.000 117.200 ;
        RECT 29.700 115.600 34.600 115.700 ;
        RECT 31.700 115.500 34.600 115.600 ;
        RECT 31.800 115.400 34.600 115.500 ;
        RECT 26.300 114.900 26.700 115.000 ;
        RECT 26.300 114.600 28.200 114.900 ;
        RECT 28.600 114.800 29.000 115.200 ;
        RECT 31.000 115.100 31.400 115.200 ;
        RECT 31.000 114.800 33.500 115.100 ;
        RECT 27.800 114.500 28.200 114.600 ;
        RECT 28.700 114.200 29.000 114.800 ;
        RECT 31.800 114.700 32.200 114.800 ;
        RECT 33.100 114.700 33.500 114.800 ;
        RECT 35.800 114.400 36.200 115.200 ;
        RECT 32.300 114.200 32.700 114.300 ;
        RECT 36.500 114.200 36.800 115.900 ;
        RECT 37.400 115.800 37.800 115.900 ;
        RECT 38.300 115.200 38.600 115.900 ;
        RECT 40.200 115.200 40.600 115.400 ;
        RECT 38.200 114.900 39.400 115.200 ;
        RECT 40.200 114.900 41.000 115.200 ;
        RECT 38.200 114.800 38.600 114.900 ;
        RECT 28.700 113.900 34.200 114.200 ;
        RECT 28.900 113.800 29.300 113.900 ;
        RECT 25.400 113.300 27.300 113.600 ;
        RECT 25.400 111.100 25.800 113.300 ;
        RECT 26.900 113.200 27.300 113.300 ;
        RECT 31.800 112.800 32.100 113.900 ;
        RECT 33.400 113.800 34.200 113.900 ;
        RECT 35.000 114.100 35.400 114.200 ;
        RECT 35.000 113.800 35.800 114.100 ;
        RECT 36.500 113.800 37.800 114.200 ;
        RECT 35.400 113.600 35.800 113.800 ;
        RECT 30.900 112.700 31.300 112.800 ;
        RECT 27.800 112.100 28.200 112.500 ;
        RECT 29.900 112.400 31.300 112.700 ;
        RECT 31.800 112.400 32.200 112.800 ;
        RECT 29.900 112.100 30.200 112.400 ;
        RECT 32.600 112.100 33.000 112.500 ;
        RECT 27.500 111.800 28.200 112.100 ;
        RECT 27.500 111.100 28.100 111.800 ;
        RECT 29.800 111.100 30.200 112.100 ;
        RECT 32.000 111.800 33.000 112.100 ;
        RECT 32.000 111.100 32.400 111.800 ;
        RECT 34.200 111.100 34.600 113.500 ;
        RECT 35.100 113.100 36.900 113.300 ;
        RECT 37.400 113.100 37.700 113.800 ;
        RECT 39.100 113.200 39.400 114.900 ;
        RECT 40.600 114.800 41.000 114.900 ;
        RECT 39.800 113.800 40.200 114.600 ;
        RECT 42.300 114.200 42.600 115.900 ;
        RECT 43.800 115.800 44.200 116.200 ;
        RECT 43.000 114.800 43.400 115.600 ;
        RECT 42.200 113.800 42.600 114.200 ;
        RECT 43.900 114.200 44.200 115.800 ;
        RECT 46.200 116.100 46.600 116.200 ;
        RECT 47.800 116.100 48.200 116.200 ;
        RECT 46.200 115.800 48.200 116.100 ;
        RECT 48.600 115.800 49.000 116.200 ;
        RECT 46.200 115.400 46.600 115.800 ;
        RECT 45.000 114.800 45.800 115.200 ;
        RECT 48.700 114.200 49.000 115.800 ;
        RECT 51.000 115.400 51.400 116.200 ;
        RECT 51.800 115.800 52.200 116.200 ;
        RECT 49.800 114.800 50.600 115.200 ;
        RECT 51.900 114.200 52.200 115.800 ;
        RECT 54.200 115.400 54.600 116.200 ;
        RECT 55.000 116.100 55.400 119.900 ;
        RECT 55.800 116.100 56.200 116.200 ;
        RECT 55.000 115.800 56.200 116.100 ;
        RECT 56.600 115.800 57.000 116.600 ;
        RECT 53.000 114.800 53.800 115.200 ;
        RECT 43.900 114.100 44.700 114.200 ;
        RECT 48.700 114.100 49.500 114.200 ;
        RECT 51.900 114.100 52.700 114.200 ;
        RECT 43.900 113.900 44.800 114.100 ;
        RECT 48.700 113.900 49.600 114.100 ;
        RECT 51.900 113.900 52.800 114.100 ;
        RECT 38.200 113.100 38.600 113.200 ;
        RECT 35.000 113.000 37.000 113.100 ;
        RECT 35.000 111.100 35.400 113.000 ;
        RECT 36.600 111.100 37.000 113.000 ;
        RECT 37.400 112.800 38.600 113.100 ;
        RECT 37.400 111.100 37.800 112.800 ;
        RECT 38.300 112.400 38.700 112.800 ;
        RECT 39.000 111.100 39.400 113.200 ;
        RECT 41.400 112.400 41.800 113.200 ;
        RECT 42.300 112.100 42.600 113.800 ;
        RECT 42.200 111.100 42.600 112.100 ;
        RECT 44.400 111.100 44.800 113.900 ;
        RECT 49.200 111.100 49.600 113.900 ;
        RECT 52.400 111.100 52.800 113.900 ;
        RECT 55.000 111.100 55.400 115.800 ;
        RECT 55.800 113.100 56.200 113.200 ;
        RECT 57.400 113.100 57.800 119.900 ;
        RECT 59.400 116.800 59.800 117.200 ;
        RECT 59.400 116.200 59.700 116.800 ;
        RECT 60.100 116.200 60.500 119.900 ;
        RECT 59.000 115.900 59.700 116.200 ;
        RECT 60.000 115.900 60.500 116.200 ;
        RECT 62.200 116.100 62.600 119.900 ;
        RECT 63.000 116.100 63.400 116.200 ;
        RECT 59.000 115.800 59.400 115.900 ;
        RECT 59.000 115.100 59.400 115.200 ;
        RECT 60.000 115.100 60.300 115.900 ;
        RECT 62.200 115.800 63.400 116.100 ;
        RECT 63.800 115.900 64.200 119.900 ;
        RECT 65.400 117.900 65.800 119.900 ;
        RECT 59.000 114.800 60.300 115.100 ;
        RECT 60.000 114.200 60.300 114.800 ;
        RECT 60.600 114.400 61.000 115.200 ;
        RECT 58.200 113.400 58.600 114.200 ;
        RECT 59.000 113.800 60.300 114.200 ;
        RECT 61.400 114.100 61.800 114.200 ;
        RECT 61.000 113.800 61.800 114.100 ;
        RECT 59.100 113.100 59.400 113.800 ;
        RECT 61.000 113.600 61.400 113.800 ;
        RECT 59.900 113.100 61.700 113.300 ;
        RECT 55.800 112.800 57.800 113.100 ;
        RECT 55.800 112.400 56.200 112.800 ;
        RECT 56.900 111.100 57.300 112.800 ;
        RECT 59.000 111.100 59.400 113.100 ;
        RECT 59.800 113.000 61.800 113.100 ;
        RECT 59.800 111.100 60.200 113.000 ;
        RECT 61.400 111.100 61.800 113.000 ;
        RECT 62.200 111.100 62.600 115.800 ;
        RECT 63.800 115.200 64.100 115.900 ;
        RECT 65.400 115.800 65.700 117.900 ;
        RECT 68.300 116.300 68.700 119.900 ;
        RECT 67.800 115.900 68.700 116.300 ;
        RECT 64.500 115.500 65.700 115.800 ;
        RECT 63.800 114.800 64.200 115.200 ;
        RECT 63.000 112.400 63.400 113.200 ;
        RECT 63.800 113.100 64.100 114.800 ;
        RECT 64.500 113.800 64.800 115.500 ;
        RECT 65.400 114.800 65.800 115.200 ;
        RECT 65.400 114.400 65.700 114.800 ;
        RECT 65.200 114.100 65.700 114.400 ;
        RECT 66.200 114.100 66.600 114.600 ;
        RECT 67.900 114.200 68.200 115.900 ;
        RECT 69.400 115.600 69.800 119.900 ;
        RECT 71.500 117.900 72.100 119.900 ;
        RECT 73.800 117.900 74.200 119.900 ;
        RECT 76.000 118.200 76.400 119.900 ;
        RECT 76.000 117.900 77.000 118.200 ;
        RECT 71.800 117.500 72.200 117.900 ;
        RECT 73.900 117.600 74.200 117.900 ;
        RECT 73.500 117.300 75.300 117.600 ;
        RECT 76.600 117.500 77.000 117.900 ;
        RECT 73.500 117.200 73.900 117.300 ;
        RECT 74.900 117.200 75.300 117.300 ;
        RECT 71.400 116.600 72.100 117.000 ;
        RECT 71.800 116.100 72.100 116.600 ;
        RECT 72.900 116.500 74.000 116.800 ;
        RECT 72.900 116.400 73.300 116.500 ;
        RECT 71.800 115.800 73.000 116.100 ;
        RECT 68.600 114.800 69.000 115.600 ;
        RECT 69.400 115.300 71.500 115.600 ;
        RECT 65.200 114.000 65.600 114.100 ;
        RECT 66.200 113.800 67.300 114.100 ;
        RECT 67.800 113.800 68.200 114.200 ;
        RECT 64.400 113.700 64.800 113.800 ;
        RECT 64.400 113.500 65.900 113.700 ;
        RECT 64.400 113.400 66.500 113.500 ;
        RECT 65.600 113.200 66.500 113.400 ;
        RECT 66.200 113.100 66.500 113.200 ;
        RECT 67.000 113.200 67.300 113.800 ;
        RECT 63.800 112.600 64.500 113.100 ;
        RECT 64.100 112.200 64.500 112.600 ;
        RECT 63.800 111.800 64.500 112.200 ;
        RECT 64.100 111.100 64.500 111.800 ;
        RECT 66.200 111.100 66.600 113.100 ;
        RECT 67.000 112.400 67.400 113.200 ;
        RECT 67.900 112.200 68.200 113.800 ;
        RECT 69.400 113.600 69.800 115.300 ;
        RECT 71.100 115.200 71.500 115.300 ;
        RECT 70.300 114.900 70.700 115.000 ;
        RECT 70.300 114.600 72.200 114.900 ;
        RECT 71.800 114.500 72.200 114.600 ;
        RECT 72.700 114.200 73.000 115.800 ;
        RECT 73.700 115.900 74.000 116.500 ;
        RECT 74.300 116.500 74.700 116.600 ;
        RECT 76.600 116.500 77.000 116.600 ;
        RECT 74.300 116.200 77.000 116.500 ;
        RECT 73.700 115.700 76.100 115.900 ;
        RECT 78.200 115.700 78.600 119.900 ;
        RECT 73.700 115.600 78.600 115.700 ;
        RECT 75.700 115.500 78.600 115.600 ;
        RECT 75.800 115.400 78.600 115.500 ;
        RECT 75.000 115.100 75.400 115.200 ;
        RECT 75.000 114.800 77.500 115.100 ;
        RECT 75.800 114.700 76.200 114.800 ;
        RECT 77.100 114.700 77.500 114.800 ;
        RECT 76.300 114.200 76.700 114.300 ;
        RECT 72.700 113.900 78.200 114.200 ;
        RECT 72.900 113.800 73.300 113.900 ;
        RECT 69.400 113.300 71.300 113.600 ;
        RECT 68.600 113.100 69.000 113.200 ;
        RECT 69.400 113.100 69.800 113.300 ;
        RECT 70.900 113.200 71.300 113.300 ;
        RECT 68.600 112.800 69.800 113.100 ;
        RECT 75.800 112.800 76.100 113.900 ;
        RECT 77.400 113.800 78.200 113.900 ;
        RECT 79.000 114.100 79.400 119.900 ;
        RECT 81.900 116.200 82.300 119.900 ;
        RECT 82.600 116.800 83.000 117.200 ;
        RECT 82.700 116.200 83.000 116.800 ;
        RECT 81.900 115.900 82.400 116.200 ;
        RECT 82.700 115.900 83.400 116.200 ;
        RECT 81.400 114.400 81.800 115.200 ;
        RECT 82.100 114.200 82.400 115.900 ;
        RECT 83.000 115.800 83.400 115.900 ;
        RECT 83.800 115.800 84.200 116.600 ;
        RECT 83.000 115.100 83.300 115.800 ;
        RECT 84.600 115.100 85.000 119.900 ;
        RECT 86.200 117.500 86.600 119.500 ;
        RECT 86.200 115.800 86.500 117.500 ;
        RECT 88.300 116.400 88.700 119.900 ;
        RECT 88.300 116.100 89.100 116.400 ;
        RECT 86.200 115.500 88.100 115.800 ;
        RECT 83.000 114.800 85.000 115.100 ;
        RECT 80.600 114.100 81.000 114.200 ;
        RECT 79.000 113.800 81.400 114.100 ;
        RECT 82.100 113.800 83.400 114.200 ;
        RECT 67.800 111.100 68.200 112.200 ;
        RECT 69.400 111.100 69.800 112.800 ;
        RECT 74.900 112.700 75.300 112.800 ;
        RECT 71.800 112.100 72.200 112.500 ;
        RECT 73.900 112.400 75.300 112.700 ;
        RECT 75.800 112.400 76.200 112.800 ;
        RECT 73.900 112.100 74.200 112.400 ;
        RECT 76.600 112.100 77.000 112.500 ;
        RECT 71.500 111.800 72.200 112.100 ;
        RECT 71.500 111.100 72.100 111.800 ;
        RECT 73.800 111.100 74.200 112.100 ;
        RECT 76.000 111.800 77.000 112.100 ;
        RECT 76.000 111.100 76.400 111.800 ;
        RECT 78.200 111.100 78.600 113.500 ;
        RECT 79.000 111.100 79.400 113.800 ;
        RECT 81.000 113.600 81.400 113.800 ;
        RECT 79.800 112.400 80.200 113.200 ;
        RECT 80.700 113.100 82.500 113.300 ;
        RECT 83.000 113.100 83.300 113.800 ;
        RECT 84.600 113.100 85.000 114.800 ;
        RECT 86.200 114.400 86.600 115.200 ;
        RECT 87.000 114.400 87.400 115.200 ;
        RECT 87.800 114.500 88.100 115.500 ;
        RECT 85.400 113.400 85.800 114.200 ;
        RECT 87.800 114.100 88.500 114.500 ;
        RECT 88.800 114.200 89.100 116.100 ;
        RECT 91.300 116.300 91.700 119.900 ;
        RECT 91.300 115.900 92.200 116.300 ;
        RECT 89.400 114.800 89.800 115.600 ;
        RECT 91.000 114.800 91.400 115.600 ;
        RECT 88.800 114.100 89.800 114.200 ;
        RECT 91.000 114.100 91.300 114.800 ;
        RECT 87.800 113.900 88.300 114.100 ;
        RECT 86.200 113.600 88.300 113.900 ;
        RECT 88.800 113.800 91.300 114.100 ;
        RECT 91.800 114.200 92.100 115.900 ;
        RECT 95.000 115.600 95.400 119.900 ;
        RECT 97.100 117.900 97.700 119.900 ;
        RECT 99.400 117.900 99.800 119.900 ;
        RECT 101.600 118.200 102.000 119.900 ;
        RECT 101.600 117.900 102.600 118.200 ;
        RECT 97.400 117.500 97.800 117.900 ;
        RECT 99.500 117.600 99.800 117.900 ;
        RECT 99.100 117.300 100.900 117.600 ;
        RECT 102.200 117.500 102.600 117.900 ;
        RECT 99.100 117.200 99.500 117.300 ;
        RECT 100.500 117.200 100.900 117.300 ;
        RECT 97.000 116.600 97.700 117.000 ;
        RECT 97.400 116.100 97.700 116.600 ;
        RECT 98.500 116.500 99.600 116.800 ;
        RECT 98.500 116.400 98.900 116.500 ;
        RECT 97.400 115.800 98.600 116.100 ;
        RECT 95.000 115.300 97.100 115.600 ;
        RECT 91.800 113.800 92.200 114.200 ;
        RECT 80.600 113.000 82.600 113.100 ;
        RECT 80.600 111.100 81.000 113.000 ;
        RECT 82.200 111.100 82.600 113.000 ;
        RECT 83.000 111.100 83.400 113.100 ;
        RECT 84.100 112.800 85.000 113.100 ;
        RECT 84.100 111.100 84.500 112.800 ;
        RECT 86.200 112.500 86.500 113.600 ;
        RECT 88.800 113.500 89.100 113.800 ;
        RECT 88.700 113.300 89.100 113.500 ;
        RECT 88.300 113.000 89.100 113.300 ;
        RECT 86.200 111.500 86.600 112.500 ;
        RECT 88.300 111.500 88.700 113.000 ;
        RECT 91.800 112.200 92.100 113.800 ;
        RECT 95.000 113.600 95.400 115.300 ;
        RECT 96.700 115.200 97.100 115.300 ;
        RECT 95.900 114.900 96.300 115.000 ;
        RECT 95.900 114.600 97.800 114.900 ;
        RECT 97.400 114.500 97.800 114.600 ;
        RECT 98.300 114.200 98.600 115.800 ;
        RECT 99.300 115.900 99.600 116.500 ;
        RECT 99.900 116.500 100.300 116.600 ;
        RECT 102.200 116.500 102.600 116.600 ;
        RECT 99.900 116.200 102.600 116.500 ;
        RECT 99.300 115.700 101.700 115.900 ;
        RECT 103.800 115.700 104.200 119.900 ;
        RECT 99.300 115.600 104.200 115.700 ;
        RECT 101.300 115.500 104.200 115.600 ;
        RECT 101.400 115.400 104.200 115.500 ;
        RECT 104.600 115.700 105.000 119.900 ;
        RECT 106.800 118.200 107.200 119.900 ;
        RECT 106.200 117.900 107.200 118.200 ;
        RECT 109.000 117.900 109.400 119.900 ;
        RECT 111.100 117.900 111.700 119.900 ;
        RECT 113.400 119.100 113.800 119.900 ;
        RECT 114.200 119.100 114.600 119.900 ;
        RECT 113.400 118.800 114.600 119.100 ;
        RECT 106.200 117.500 106.600 117.900 ;
        RECT 109.000 117.600 109.300 117.900 ;
        RECT 107.900 117.300 109.700 117.600 ;
        RECT 111.000 117.500 111.400 117.900 ;
        RECT 107.900 117.200 108.300 117.300 ;
        RECT 109.300 117.200 109.700 117.300 ;
        RECT 106.200 116.500 106.600 116.600 ;
        RECT 108.500 116.500 108.900 116.600 ;
        RECT 106.200 116.200 108.900 116.500 ;
        RECT 109.200 116.500 110.300 116.800 ;
        RECT 109.200 115.900 109.500 116.500 ;
        RECT 109.900 116.400 110.300 116.500 ;
        RECT 111.100 116.600 111.800 117.000 ;
        RECT 111.100 116.100 111.400 116.600 ;
        RECT 107.100 115.700 109.500 115.900 ;
        RECT 104.600 115.600 109.500 115.700 ;
        RECT 110.200 115.800 111.400 116.100 ;
        RECT 104.600 115.500 107.500 115.600 ;
        RECT 104.600 115.400 107.400 115.500 ;
        RECT 110.200 115.200 110.500 115.800 ;
        RECT 113.400 115.600 113.800 118.800 ;
        RECT 111.700 115.300 113.800 115.600 ;
        RECT 111.700 115.200 112.100 115.300 ;
        RECT 100.600 115.100 101.000 115.200 ;
        RECT 107.800 115.100 108.200 115.200 ;
        RECT 100.600 114.800 103.100 115.100 ;
        RECT 101.400 114.700 101.800 114.800 ;
        RECT 102.700 114.700 103.100 114.800 ;
        RECT 105.700 114.800 108.200 115.100 ;
        RECT 110.200 114.800 110.600 115.200 ;
        RECT 112.500 114.900 112.900 115.000 ;
        RECT 105.700 114.700 106.100 114.800 ;
        RECT 101.900 114.200 102.300 114.300 ;
        RECT 106.500 114.200 106.900 114.300 ;
        RECT 110.200 114.200 110.500 114.800 ;
        RECT 111.000 114.600 112.900 114.900 ;
        RECT 111.000 114.500 111.400 114.600 ;
        RECT 98.200 114.100 103.800 114.200 ;
        RECT 105.000 114.100 110.500 114.200 ;
        RECT 98.200 113.900 110.500 114.100 ;
        RECT 98.200 113.800 98.900 113.900 ;
        RECT 95.000 113.300 96.900 113.600 ;
        RECT 92.600 112.400 93.000 113.200 ;
        RECT 91.800 111.100 92.200 112.200 ;
        RECT 95.000 111.100 95.400 113.300 ;
        RECT 96.500 113.200 96.900 113.300 ;
        RECT 101.400 112.800 101.700 113.900 ;
        RECT 103.000 113.800 105.800 113.900 ;
        RECT 100.500 112.700 100.900 112.800 ;
        RECT 97.400 112.100 97.800 112.500 ;
        RECT 99.500 112.400 100.900 112.700 ;
        RECT 101.400 112.400 101.800 112.800 ;
        RECT 99.500 112.100 99.800 112.400 ;
        RECT 102.200 112.100 102.600 112.500 ;
        RECT 97.100 111.800 97.800 112.100 ;
        RECT 97.100 111.100 97.700 111.800 ;
        RECT 99.400 111.100 99.800 112.100 ;
        RECT 101.600 111.800 102.600 112.100 ;
        RECT 101.600 111.100 102.000 111.800 ;
        RECT 103.800 111.100 104.200 113.500 ;
        RECT 104.600 111.100 105.000 113.500 ;
        RECT 107.100 112.800 107.400 113.900 ;
        RECT 109.900 113.800 110.300 113.900 ;
        RECT 113.400 113.600 113.800 115.300 ;
        RECT 111.900 113.300 113.800 113.600 ;
        RECT 111.900 113.200 112.300 113.300 ;
        RECT 106.200 112.100 106.600 112.500 ;
        RECT 107.000 112.400 107.400 112.800 ;
        RECT 107.900 112.700 108.300 112.800 ;
        RECT 107.900 112.400 109.300 112.700 ;
        RECT 109.000 112.100 109.300 112.400 ;
        RECT 111.000 112.100 111.400 112.500 ;
        RECT 106.200 111.800 107.200 112.100 ;
        RECT 106.800 111.100 107.200 111.800 ;
        RECT 109.000 111.100 109.400 112.100 ;
        RECT 111.000 111.800 111.700 112.100 ;
        RECT 111.100 111.100 111.700 111.800 ;
        RECT 113.400 111.100 113.800 113.300 ;
        RECT 114.200 115.600 114.600 118.800 ;
        RECT 116.300 117.900 116.900 119.900 ;
        RECT 118.600 117.900 119.000 119.900 ;
        RECT 120.800 118.200 121.200 119.900 ;
        RECT 120.800 117.900 121.800 118.200 ;
        RECT 116.600 117.500 117.000 117.900 ;
        RECT 118.700 117.600 119.000 117.900 ;
        RECT 118.300 117.300 120.100 117.600 ;
        RECT 121.400 117.500 121.800 117.900 ;
        RECT 118.300 117.200 118.700 117.300 ;
        RECT 119.700 117.200 120.100 117.300 ;
        RECT 116.200 116.600 116.900 117.000 ;
        RECT 116.600 116.100 116.900 116.600 ;
        RECT 117.700 116.500 118.800 116.800 ;
        RECT 117.700 116.400 118.100 116.500 ;
        RECT 116.600 115.800 117.800 116.100 ;
        RECT 114.200 115.300 116.300 115.600 ;
        RECT 114.200 113.600 114.600 115.300 ;
        RECT 115.900 115.200 116.300 115.300 ;
        RECT 117.500 115.200 117.800 115.800 ;
        RECT 118.500 115.900 118.800 116.500 ;
        RECT 119.100 116.500 119.500 116.600 ;
        RECT 121.400 116.500 121.800 116.600 ;
        RECT 119.100 116.200 121.800 116.500 ;
        RECT 118.500 115.700 120.900 115.900 ;
        RECT 123.000 115.700 123.400 119.900 ;
        RECT 125.100 116.300 125.500 119.900 ;
        RECT 128.100 116.400 128.500 119.900 ;
        RECT 130.200 117.500 130.600 119.500 ;
        RECT 124.600 115.900 125.500 116.300 ;
        RECT 127.700 116.100 128.500 116.400 ;
        RECT 118.500 115.600 123.400 115.700 ;
        RECT 120.500 115.500 123.400 115.600 ;
        RECT 120.600 115.400 123.400 115.500 ;
        RECT 115.100 114.900 115.500 115.000 ;
        RECT 115.100 114.600 117.000 114.900 ;
        RECT 117.400 114.800 117.800 115.200 ;
        RECT 119.800 115.100 120.200 115.200 ;
        RECT 119.800 114.800 122.300 115.100 ;
        RECT 116.600 114.500 117.000 114.600 ;
        RECT 117.500 114.200 117.800 114.800 ;
        RECT 120.600 114.700 121.000 114.800 ;
        RECT 121.900 114.700 122.300 114.800 ;
        RECT 121.100 114.200 121.500 114.300 ;
        RECT 124.700 114.200 125.000 115.900 ;
        RECT 127.700 115.800 128.200 116.100 ;
        RECT 130.300 115.800 130.600 117.500 ;
        RECT 131.000 115.800 131.400 116.600 ;
        RECT 125.400 114.800 125.800 115.600 ;
        RECT 126.200 115.100 126.600 115.200 ;
        RECT 127.000 115.100 127.400 115.600 ;
        RECT 126.200 114.800 127.400 115.100 ;
        RECT 127.700 114.200 128.000 115.800 ;
        RECT 128.700 115.500 130.600 115.800 ;
        RECT 128.700 114.500 129.000 115.500 ;
        RECT 117.500 113.900 123.000 114.200 ;
        RECT 117.700 113.800 118.100 113.900 ;
        RECT 114.200 113.300 116.100 113.600 ;
        RECT 114.200 111.100 114.600 113.300 ;
        RECT 115.700 113.200 116.100 113.300 ;
        RECT 120.600 112.800 120.900 113.900 ;
        RECT 122.200 113.800 123.000 113.900 ;
        RECT 124.600 114.100 125.000 114.200 ;
        RECT 125.400 114.100 125.800 114.200 ;
        RECT 124.600 113.800 125.800 114.100 ;
        RECT 127.000 113.800 128.000 114.200 ;
        RECT 128.300 114.100 129.000 114.500 ;
        RECT 129.400 114.400 129.800 115.200 ;
        RECT 130.200 114.400 130.600 115.200 ;
        RECT 119.700 112.700 120.100 112.800 ;
        RECT 116.600 112.100 117.000 112.500 ;
        RECT 118.700 112.400 120.100 112.700 ;
        RECT 120.600 112.400 121.000 112.800 ;
        RECT 118.700 112.100 119.000 112.400 ;
        RECT 121.400 112.100 121.800 112.500 ;
        RECT 116.300 111.800 117.000 112.100 ;
        RECT 116.300 111.100 116.900 111.800 ;
        RECT 118.600 111.100 119.000 112.100 ;
        RECT 120.800 111.800 121.800 112.100 ;
        RECT 120.800 111.100 121.200 111.800 ;
        RECT 123.000 111.100 123.400 113.500 ;
        RECT 123.800 112.400 124.200 113.200 ;
        RECT 124.700 112.100 125.000 113.800 ;
        RECT 127.700 113.500 128.000 113.800 ;
        RECT 128.500 113.900 129.000 114.100 ;
        RECT 128.500 113.600 130.600 113.900 ;
        RECT 127.700 113.300 128.100 113.500 ;
        RECT 127.700 113.000 128.500 113.300 ;
        RECT 124.600 111.100 125.000 112.100 ;
        RECT 128.100 111.500 128.500 113.000 ;
        RECT 130.300 112.500 130.600 113.600 ;
        RECT 131.800 113.100 132.200 119.900 ;
        RECT 134.700 116.300 135.100 119.900 ;
        RECT 134.200 115.900 135.100 116.300 ;
        RECT 134.300 114.200 134.600 115.900 ;
        RECT 135.000 114.800 135.400 115.600 ;
        RECT 136.600 115.100 137.000 119.900 ;
        RECT 138.600 116.800 139.000 117.200 ;
        RECT 137.400 115.800 137.800 116.600 ;
        RECT 138.600 116.200 138.900 116.800 ;
        RECT 139.300 116.200 139.700 119.900 ;
        RECT 138.200 115.900 138.900 116.200 ;
        RECT 139.200 115.900 139.700 116.200 ;
        RECT 138.200 115.800 138.600 115.900 ;
        RECT 138.200 115.100 138.500 115.800 ;
        RECT 136.600 114.800 138.500 115.100 ;
        RECT 132.600 114.100 133.000 114.200 ;
        RECT 134.200 114.100 134.600 114.200 ;
        RECT 132.600 113.800 134.600 114.100 ;
        RECT 132.600 113.400 133.000 113.800 ;
        RECT 130.200 111.500 130.600 112.500 ;
        RECT 131.300 112.800 132.200 113.100 ;
        RECT 131.300 112.200 131.700 112.800 ;
        RECT 133.400 112.400 133.800 113.200 ;
        RECT 131.300 111.800 132.200 112.200 ;
        RECT 134.300 112.100 134.600 113.800 ;
        RECT 135.800 113.400 136.200 114.200 ;
        RECT 136.600 113.100 137.000 114.800 ;
        RECT 139.200 114.200 139.500 115.900 ;
        RECT 139.800 114.400 140.200 115.200 ;
        RECT 138.200 113.800 139.500 114.200 ;
        RECT 140.600 114.100 141.000 114.200 ;
        RECT 141.400 114.100 141.800 119.900 ;
        RECT 140.200 113.800 141.800 114.100 ;
        RECT 138.300 113.100 138.600 113.800 ;
        RECT 140.200 113.600 140.600 113.800 ;
        RECT 139.100 113.100 140.900 113.300 ;
        RECT 136.600 112.800 137.500 113.100 ;
        RECT 131.300 111.100 131.700 111.800 ;
        RECT 134.200 111.100 134.600 112.100 ;
        RECT 137.100 111.100 137.500 112.800 ;
        RECT 138.200 111.100 138.600 113.100 ;
        RECT 139.000 113.000 141.000 113.100 ;
        RECT 139.000 111.100 139.400 113.000 ;
        RECT 140.600 111.100 141.000 113.000 ;
        RECT 141.400 111.100 141.800 113.800 ;
        RECT 142.200 112.400 142.600 113.200 ;
        RECT 143.000 111.100 143.400 119.900 ;
        RECT 146.200 115.600 146.600 119.900 ;
        RECT 148.300 117.900 148.900 119.900 ;
        RECT 150.600 117.900 151.000 119.900 ;
        RECT 152.800 118.200 153.200 119.900 ;
        RECT 152.800 117.900 153.800 118.200 ;
        RECT 148.600 117.500 149.000 117.900 ;
        RECT 150.700 117.600 151.000 117.900 ;
        RECT 150.300 117.300 152.100 117.600 ;
        RECT 153.400 117.500 153.800 117.900 ;
        RECT 150.300 117.200 150.700 117.300 ;
        RECT 151.700 117.200 152.100 117.300 ;
        RECT 148.200 116.600 148.900 117.000 ;
        RECT 148.600 116.100 148.900 116.600 ;
        RECT 149.700 116.500 150.800 116.800 ;
        RECT 149.700 116.400 150.100 116.500 ;
        RECT 148.600 115.800 149.800 116.100 ;
        RECT 146.200 115.300 148.300 115.600 ;
        RECT 146.200 113.600 146.600 115.300 ;
        RECT 147.900 115.200 148.300 115.300 ;
        RECT 147.100 114.900 147.500 115.000 ;
        RECT 147.100 114.600 149.000 114.900 ;
        RECT 148.600 114.500 149.000 114.600 ;
        RECT 149.500 114.200 149.800 115.800 ;
        RECT 150.500 115.900 150.800 116.500 ;
        RECT 151.100 116.500 151.500 116.600 ;
        RECT 153.400 116.500 153.800 116.600 ;
        RECT 151.100 116.200 153.800 116.500 ;
        RECT 150.500 115.700 152.900 115.900 ;
        RECT 155.000 115.700 155.400 119.900 ;
        RECT 156.600 117.900 157.000 119.900 ;
        RECT 150.500 115.600 155.400 115.700 ;
        RECT 152.500 115.500 155.400 115.600 ;
        RECT 156.700 115.800 157.000 117.900 ;
        RECT 158.200 115.900 158.600 119.900 ;
        RECT 156.700 115.500 157.900 115.800 ;
        RECT 152.600 115.400 155.400 115.500 ;
        RECT 151.800 115.100 152.200 115.200 ;
        RECT 151.800 114.800 154.300 115.100 ;
        RECT 156.600 114.800 157.000 115.200 ;
        RECT 152.600 114.700 153.000 114.800 ;
        RECT 153.900 114.700 154.300 114.800 ;
        RECT 153.100 114.200 153.500 114.300 ;
        RECT 149.500 113.900 155.000 114.200 ;
        RECT 149.700 113.800 150.100 113.900 ;
        RECT 146.200 113.300 148.100 113.600 ;
        RECT 143.800 113.100 144.200 113.200 ;
        RECT 145.400 113.100 145.800 113.200 ;
        RECT 143.800 112.800 145.800 113.100 ;
        RECT 143.800 112.400 144.200 112.800 ;
        RECT 146.200 111.100 146.600 113.300 ;
        RECT 147.700 113.200 148.100 113.300 ;
        RECT 152.600 112.800 152.900 113.900 ;
        RECT 154.200 113.800 155.000 113.900 ;
        RECT 155.800 113.800 156.200 114.600 ;
        RECT 156.700 114.400 157.000 114.800 ;
        RECT 156.700 114.100 157.200 114.400 ;
        RECT 156.800 114.000 157.200 114.100 ;
        RECT 157.600 113.800 157.900 115.500 ;
        RECT 158.300 115.200 158.600 115.900 ;
        RECT 158.200 114.800 158.600 115.200 ;
        RECT 157.600 113.700 158.000 113.800 ;
        RECT 156.500 113.500 158.000 113.700 ;
        RECT 151.700 112.700 152.100 112.800 ;
        RECT 148.600 112.100 149.000 112.500 ;
        RECT 150.700 112.400 152.100 112.700 ;
        RECT 152.600 112.400 153.000 112.800 ;
        RECT 150.700 112.100 151.000 112.400 ;
        RECT 153.400 112.100 153.800 112.500 ;
        RECT 148.300 111.800 149.000 112.100 ;
        RECT 148.300 111.100 148.900 111.800 ;
        RECT 150.600 111.100 151.000 112.100 ;
        RECT 152.800 111.800 153.800 112.100 ;
        RECT 152.800 111.100 153.200 111.800 ;
        RECT 155.000 111.100 155.400 113.500 ;
        RECT 155.900 113.400 158.000 113.500 ;
        RECT 155.900 113.200 156.800 113.400 ;
        RECT 155.900 113.100 156.200 113.200 ;
        RECT 158.300 113.100 158.600 114.800 ;
        RECT 155.800 111.100 156.200 113.100 ;
        RECT 157.900 112.600 158.600 113.100 ;
        RECT 159.000 115.600 159.400 119.900 ;
        RECT 161.100 117.900 161.700 119.900 ;
        RECT 163.400 117.900 163.800 119.900 ;
        RECT 165.600 118.200 166.000 119.900 ;
        RECT 165.600 117.900 166.600 118.200 ;
        RECT 161.400 117.500 161.800 117.900 ;
        RECT 163.500 117.600 163.800 117.900 ;
        RECT 163.100 117.300 164.900 117.600 ;
        RECT 166.200 117.500 166.600 117.900 ;
        RECT 163.100 117.200 163.500 117.300 ;
        RECT 164.500 117.200 164.900 117.300 ;
        RECT 161.000 116.600 161.700 117.000 ;
        RECT 161.400 116.100 161.700 116.600 ;
        RECT 162.500 116.500 163.600 116.800 ;
        RECT 162.500 116.400 162.900 116.500 ;
        RECT 161.400 115.800 162.600 116.100 ;
        RECT 159.000 115.300 161.100 115.600 ;
        RECT 159.000 113.600 159.400 115.300 ;
        RECT 160.700 115.200 161.100 115.300 ;
        RECT 159.900 114.900 160.300 115.000 ;
        RECT 159.900 114.600 161.800 114.900 ;
        RECT 161.400 114.500 161.800 114.600 ;
        RECT 162.300 114.200 162.600 115.800 ;
        RECT 163.300 115.900 163.600 116.500 ;
        RECT 163.900 116.500 164.300 116.600 ;
        RECT 166.200 116.500 166.600 116.600 ;
        RECT 163.900 116.200 166.600 116.500 ;
        RECT 163.300 115.700 165.700 115.900 ;
        RECT 167.800 115.700 168.200 119.900 ;
        RECT 163.300 115.600 168.200 115.700 ;
        RECT 165.300 115.500 168.200 115.600 ;
        RECT 165.400 115.400 168.200 115.500 ;
        RECT 168.600 115.600 169.000 119.900 ;
        RECT 170.700 117.900 171.300 119.900 ;
        RECT 173.000 117.900 173.400 119.900 ;
        RECT 175.200 118.200 175.600 119.900 ;
        RECT 175.200 117.900 176.200 118.200 ;
        RECT 171.000 117.500 171.400 117.900 ;
        RECT 173.100 117.600 173.400 117.900 ;
        RECT 172.700 117.300 174.500 117.600 ;
        RECT 175.800 117.500 176.200 117.900 ;
        RECT 172.700 117.200 173.100 117.300 ;
        RECT 174.100 117.200 174.500 117.300 ;
        RECT 170.600 116.600 171.300 117.000 ;
        RECT 171.000 116.100 171.300 116.600 ;
        RECT 172.100 116.500 173.200 116.800 ;
        RECT 172.100 116.400 172.500 116.500 ;
        RECT 171.000 115.800 172.200 116.100 ;
        RECT 168.600 115.300 170.700 115.600 ;
        RECT 164.600 115.100 165.000 115.200 ;
        RECT 164.600 114.800 167.100 115.100 ;
        RECT 165.400 114.700 165.800 114.800 ;
        RECT 166.700 114.700 167.100 114.800 ;
        RECT 165.900 114.200 166.300 114.300 ;
        RECT 162.300 113.900 167.800 114.200 ;
        RECT 162.500 113.800 162.900 113.900 ;
        RECT 159.000 113.300 160.900 113.600 ;
        RECT 157.900 112.200 158.300 112.600 ;
        RECT 157.900 111.800 158.600 112.200 ;
        RECT 157.900 111.100 158.300 111.800 ;
        RECT 159.000 111.100 159.400 113.300 ;
        RECT 160.500 113.200 160.900 113.300 ;
        RECT 165.400 112.800 165.700 113.900 ;
        RECT 167.000 113.800 167.800 113.900 ;
        RECT 168.600 113.600 169.000 115.300 ;
        RECT 170.300 115.200 170.700 115.300 ;
        RECT 169.500 114.900 169.900 115.000 ;
        RECT 169.500 114.600 171.400 114.900 ;
        RECT 171.000 114.500 171.400 114.600 ;
        RECT 171.900 114.200 172.200 115.800 ;
        RECT 172.900 115.900 173.200 116.500 ;
        RECT 173.500 116.500 173.900 116.600 ;
        RECT 175.800 116.500 176.200 116.600 ;
        RECT 173.500 116.200 176.200 116.500 ;
        RECT 172.900 115.700 175.300 115.900 ;
        RECT 177.400 115.700 177.800 119.900 ;
        RECT 180.100 116.400 180.500 119.900 ;
        RECT 182.200 117.500 182.600 119.500 ;
        RECT 172.900 115.600 177.800 115.700 ;
        RECT 179.700 116.100 180.500 116.400 ;
        RECT 179.700 115.800 180.200 116.100 ;
        RECT 182.300 115.800 182.600 117.500 ;
        RECT 183.400 116.800 183.800 117.200 ;
        RECT 183.400 116.200 183.700 116.800 ;
        RECT 184.100 116.200 184.500 119.900 ;
        RECT 183.000 115.900 183.700 116.200 ;
        RECT 184.000 115.900 184.500 116.200 ;
        RECT 186.200 116.200 186.600 119.900 ;
        RECT 188.600 116.200 189.000 119.900 ;
        RECT 190.200 116.200 190.600 119.900 ;
        RECT 186.200 115.900 187.300 116.200 ;
        RECT 188.600 115.900 190.600 116.200 ;
        RECT 191.000 115.900 191.400 119.900 ;
        RECT 191.800 116.200 192.200 119.900 ;
        RECT 191.800 115.900 192.900 116.200 ;
        RECT 193.400 115.900 193.800 119.900 ;
        RECT 183.000 115.800 183.400 115.900 ;
        RECT 174.900 115.500 177.800 115.600 ;
        RECT 175.000 115.400 177.800 115.500 ;
        RECT 174.200 115.100 174.600 115.200 ;
        RECT 174.200 114.800 176.700 115.100 ;
        RECT 179.000 114.800 179.400 115.600 ;
        RECT 175.000 114.700 175.400 114.800 ;
        RECT 176.300 114.700 176.700 114.800 ;
        RECT 175.500 114.200 175.900 114.300 ;
        RECT 179.700 114.200 180.000 115.800 ;
        RECT 180.700 115.500 182.600 115.800 ;
        RECT 180.700 114.500 181.000 115.500 ;
        RECT 184.000 115.200 184.300 115.900 ;
        RECT 187.000 115.600 187.300 115.900 ;
        RECT 187.000 115.200 187.600 115.600 ;
        RECT 189.000 115.200 189.400 115.400 ;
        RECT 191.000 115.200 191.300 115.900 ;
        RECT 192.600 115.600 192.900 115.900 ;
        RECT 192.600 115.200 193.200 115.600 ;
        RECT 171.900 113.900 177.400 114.200 ;
        RECT 172.100 113.800 172.500 113.900 ;
        RECT 164.500 112.700 164.900 112.800 ;
        RECT 161.400 112.100 161.800 112.500 ;
        RECT 163.500 112.400 164.900 112.700 ;
        RECT 165.400 112.400 165.800 112.800 ;
        RECT 163.500 112.100 163.800 112.400 ;
        RECT 166.200 112.100 166.600 112.500 ;
        RECT 161.100 111.800 161.800 112.100 ;
        RECT 161.100 111.100 161.700 111.800 ;
        RECT 163.400 111.100 163.800 112.100 ;
        RECT 165.600 111.800 166.600 112.100 ;
        RECT 165.600 111.100 166.000 111.800 ;
        RECT 167.800 111.100 168.200 113.500 ;
        RECT 168.600 113.300 170.500 113.600 ;
        RECT 168.600 111.100 169.000 113.300 ;
        RECT 170.100 113.200 170.500 113.300 ;
        RECT 175.000 112.800 175.300 113.900 ;
        RECT 176.600 113.800 177.400 113.900 ;
        RECT 179.000 113.800 180.000 114.200 ;
        RECT 180.300 114.100 181.000 114.500 ;
        RECT 181.400 114.400 181.800 115.200 ;
        RECT 182.200 114.400 182.600 115.200 ;
        RECT 183.800 114.800 184.300 115.200 ;
        RECT 184.000 114.200 184.300 114.800 ;
        RECT 184.600 114.400 185.000 115.200 ;
        RECT 186.200 114.400 186.600 115.200 ;
        RECT 179.700 113.500 180.000 113.800 ;
        RECT 180.500 113.900 181.000 114.100 ;
        RECT 180.500 113.600 182.600 113.900 ;
        RECT 183.000 113.800 184.300 114.200 ;
        RECT 185.400 114.100 185.800 114.200 ;
        RECT 185.000 113.800 185.800 114.100 ;
        RECT 174.100 112.700 174.500 112.800 ;
        RECT 171.000 112.100 171.400 112.500 ;
        RECT 173.100 112.400 174.500 112.700 ;
        RECT 175.000 112.400 175.400 112.800 ;
        RECT 173.100 112.100 173.400 112.400 ;
        RECT 175.800 112.100 176.200 112.500 ;
        RECT 170.700 111.800 171.400 112.100 ;
        RECT 170.700 111.100 171.300 111.800 ;
        RECT 173.000 111.100 173.400 112.100 ;
        RECT 175.200 111.800 176.200 112.100 ;
        RECT 175.200 111.100 175.600 111.800 ;
        RECT 177.400 111.100 177.800 113.500 ;
        RECT 179.700 113.300 180.100 113.500 ;
        RECT 179.700 113.000 180.500 113.300 ;
        RECT 180.100 111.500 180.500 113.000 ;
        RECT 182.300 112.500 182.600 113.600 ;
        RECT 183.100 113.100 183.400 113.800 ;
        RECT 185.000 113.600 185.400 113.800 ;
        RECT 187.000 113.700 187.300 115.200 ;
        RECT 188.600 114.900 189.400 115.200 ;
        RECT 190.200 114.900 191.400 115.200 ;
        RECT 188.600 114.800 189.000 114.900 ;
        RECT 190.200 114.800 190.600 114.900 ;
        RECT 191.000 114.800 191.400 114.900 ;
        RECT 189.400 113.800 189.800 114.600 ;
        RECT 186.200 113.400 187.300 113.700 ;
        RECT 183.900 113.100 185.700 113.300 ;
        RECT 182.200 111.500 182.600 112.500 ;
        RECT 183.000 111.100 183.400 113.100 ;
        RECT 183.800 113.000 185.800 113.100 ;
        RECT 183.800 111.100 184.200 113.000 ;
        RECT 185.400 111.100 185.800 113.000 ;
        RECT 186.200 111.100 186.600 113.400 ;
        RECT 190.200 113.100 190.500 114.800 ;
        RECT 192.600 113.700 192.900 115.200 ;
        RECT 193.500 114.800 193.800 115.900 ;
        RECT 191.800 113.400 192.900 113.700 ;
        RECT 190.200 111.100 190.600 113.100 ;
        RECT 191.000 112.800 191.400 113.200 ;
        RECT 190.900 112.400 191.300 112.800 ;
        RECT 191.800 111.100 192.200 113.400 ;
        RECT 193.400 111.100 193.800 114.800 ;
        RECT 1.900 108.200 2.300 109.900 ;
        RECT 1.400 107.900 2.300 108.200 ;
        RECT 3.000 107.900 3.400 109.900 ;
        RECT 3.800 108.000 4.200 109.900 ;
        RECT 5.400 108.000 5.800 109.900 ;
        RECT 3.800 107.900 5.800 108.000 ;
        RECT 0.600 106.800 1.000 107.600 ;
        RECT 1.400 106.100 1.800 107.900 ;
        RECT 3.100 107.200 3.400 107.900 ;
        RECT 3.900 107.700 5.700 107.900 ;
        RECT 5.000 107.200 5.400 107.400 ;
        RECT 3.000 106.800 4.300 107.200 ;
        RECT 5.000 107.100 5.800 107.200 ;
        RECT 6.200 107.100 6.600 109.900 ;
        RECT 7.000 107.800 7.400 108.600 ;
        RECT 7.800 107.900 8.200 109.900 ;
        RECT 9.900 108.400 10.300 109.900 ;
        RECT 11.800 108.900 12.200 109.900 ;
        RECT 9.900 107.900 10.600 108.400 ;
        RECT 7.900 107.800 8.200 107.900 ;
        RECT 7.900 107.600 8.800 107.800 ;
        RECT 7.900 107.500 10.000 107.600 ;
        RECT 8.500 107.300 10.000 107.500 ;
        RECT 9.600 107.200 10.000 107.300 ;
        RECT 5.000 106.900 6.600 107.100 ;
        RECT 5.400 106.800 6.600 106.900 ;
        RECT 1.400 105.800 3.300 106.100 ;
        RECT 1.400 101.100 1.800 105.800 ;
        RECT 3.000 105.200 3.300 105.800 ;
        RECT 2.200 104.400 2.600 105.200 ;
        RECT 3.000 105.100 3.400 105.200 ;
        RECT 4.000 105.100 4.300 106.800 ;
        RECT 4.600 106.100 5.000 106.600 ;
        RECT 5.400 106.100 5.800 106.200 ;
        RECT 4.600 105.800 5.800 106.100 ;
        RECT 3.000 104.800 3.700 105.100 ;
        RECT 4.000 104.800 4.500 105.100 ;
        RECT 3.400 104.200 3.700 104.800 ;
        RECT 3.400 103.800 3.800 104.200 ;
        RECT 4.100 101.100 4.500 104.800 ;
        RECT 6.200 101.100 6.600 106.800 ;
        RECT 7.800 106.400 8.200 107.200 ;
        RECT 8.600 106.600 9.200 107.000 ;
        RECT 8.700 106.200 9.000 106.600 ;
        RECT 8.600 105.800 9.000 106.200 ;
        RECT 9.600 105.500 9.900 107.200 ;
        RECT 10.300 106.200 10.600 107.900 ;
        RECT 11.000 107.800 11.400 108.600 ;
        RECT 11.900 107.200 12.200 108.900 ;
        RECT 13.400 109.600 15.400 109.900 ;
        RECT 13.400 107.900 13.800 109.600 ;
        RECT 14.200 107.900 14.600 109.300 ;
        RECT 15.000 108.000 15.400 109.600 ;
        RECT 16.600 108.000 17.000 109.900 ;
        RECT 18.700 108.200 19.100 109.900 ;
        RECT 15.000 107.900 17.000 108.000 ;
        RECT 18.200 107.900 19.100 108.200 ;
        RECT 19.800 107.900 20.200 109.900 ;
        RECT 20.600 108.000 21.000 109.900 ;
        RECT 22.200 108.000 22.600 109.900 ;
        RECT 20.600 107.900 22.600 108.000 ;
        RECT 14.200 107.200 14.500 107.900 ;
        RECT 15.100 107.700 16.900 107.900 ;
        RECT 16.200 107.200 16.600 107.400 ;
        RECT 11.800 106.800 12.200 107.200 ;
        RECT 10.200 106.100 10.600 106.200 ;
        RECT 11.000 106.100 11.400 106.200 ;
        RECT 10.200 105.800 11.400 106.100 ;
        RECT 8.700 105.200 9.900 105.500 ;
        RECT 8.700 103.100 9.000 105.200 ;
        RECT 10.300 105.100 10.600 105.800 ;
        RECT 11.900 105.100 12.200 106.800 ;
        RECT 13.400 106.400 13.800 107.200 ;
        RECT 14.200 106.900 15.400 107.200 ;
        RECT 16.200 106.900 17.000 107.200 ;
        RECT 15.000 106.800 15.400 106.900 ;
        RECT 16.600 106.800 17.000 106.900 ;
        RECT 17.400 106.800 17.800 107.600 ;
        RECT 12.600 105.400 13.000 106.200 ;
        RECT 14.200 105.800 14.600 106.600 ;
        RECT 15.100 105.100 15.400 106.800 ;
        RECT 15.800 105.800 16.200 106.600 ;
        RECT 18.200 106.100 18.600 107.900 ;
        RECT 19.900 107.200 20.200 107.900 ;
        RECT 20.700 107.700 22.500 107.900 ;
        RECT 21.800 107.200 22.200 107.400 ;
        RECT 19.800 106.800 21.100 107.200 ;
        RECT 21.800 107.100 22.600 107.200 ;
        RECT 23.000 107.100 23.400 109.900 ;
        RECT 23.800 107.800 24.200 108.600 ;
        RECT 24.600 107.900 25.000 109.900 ;
        RECT 26.800 108.100 27.600 109.900 ;
        RECT 24.600 107.600 25.900 107.900 ;
        RECT 25.500 107.500 25.900 107.600 ;
        RECT 26.200 107.400 27.000 107.800 ;
        RECT 21.800 106.900 23.400 107.100 ;
        RECT 22.200 106.800 23.400 106.900 ;
        RECT 23.800 107.100 24.200 107.200 ;
        RECT 24.600 107.100 25.400 107.200 ;
        RECT 27.300 107.100 27.600 108.100 ;
        RECT 29.400 107.900 29.800 109.900 ;
        RECT 31.500 108.200 31.900 109.900 ;
        RECT 27.900 107.400 28.300 107.800 ;
        RECT 28.600 107.600 29.800 107.900 ;
        RECT 31.000 107.900 31.900 108.200 ;
        RECT 32.600 107.900 33.000 109.900 ;
        RECT 33.400 108.000 33.800 109.900 ;
        RECT 35.000 108.000 35.400 109.900 ;
        RECT 33.400 107.900 35.400 108.000 ;
        RECT 28.600 107.500 29.000 107.600 ;
        RECT 23.800 107.000 25.700 107.100 ;
        RECT 23.800 106.800 26.800 107.000 ;
        RECT 18.200 105.800 20.100 106.100 ;
        RECT 8.600 101.100 9.000 103.100 ;
        RECT 10.200 101.100 10.600 105.100 ;
        RECT 11.800 104.700 12.700 105.100 ;
        RECT 12.300 104.200 12.700 104.700 ;
        RECT 12.300 103.800 13.000 104.200 ;
        RECT 12.300 101.100 12.700 103.800 ;
        RECT 14.700 102.200 15.700 105.100 ;
        RECT 14.700 101.800 16.200 102.200 ;
        RECT 14.700 101.100 15.700 101.800 ;
        RECT 18.200 101.100 18.600 105.800 ;
        RECT 19.800 105.200 20.100 105.800 ;
        RECT 19.000 104.400 19.400 105.200 ;
        RECT 19.800 105.100 20.200 105.200 ;
        RECT 20.800 105.100 21.100 106.800 ;
        RECT 21.400 106.100 21.800 106.600 ;
        RECT 22.200 106.100 22.600 106.200 ;
        RECT 21.400 105.800 22.600 106.100 ;
        RECT 19.800 104.800 20.500 105.100 ;
        RECT 20.800 104.800 21.300 105.100 ;
        RECT 20.200 104.200 20.500 104.800 ;
        RECT 20.200 103.800 20.600 104.200 ;
        RECT 20.900 101.100 21.300 104.800 ;
        RECT 23.000 101.100 23.400 106.800 ;
        RECT 25.400 106.700 26.800 106.800 ;
        RECT 26.400 106.600 26.800 106.700 ;
        RECT 27.100 106.800 27.600 107.100 ;
        RECT 28.000 107.200 28.300 107.400 ;
        RECT 28.000 106.800 28.400 107.200 ;
        RECT 29.000 106.800 29.800 107.200 ;
        RECT 30.200 106.800 30.600 107.600 ;
        RECT 27.100 106.200 27.400 106.800 ;
        RECT 25.700 106.100 26.100 106.200 ;
        RECT 25.700 105.800 26.500 106.100 ;
        RECT 27.000 105.800 27.400 106.200 ;
        RECT 26.100 105.700 26.500 105.800 ;
        RECT 27.100 105.100 27.400 105.800 ;
        RECT 31.000 106.100 31.400 107.900 ;
        RECT 32.700 107.200 33.000 107.900 ;
        RECT 33.500 107.700 35.300 107.900 ;
        RECT 34.600 107.200 35.000 107.400 ;
        RECT 32.600 106.800 33.900 107.200 ;
        RECT 34.600 107.100 35.400 107.200 ;
        RECT 35.800 107.100 36.200 109.900 ;
        RECT 36.600 107.800 37.000 108.600 ;
        RECT 38.700 108.200 39.100 109.900 ;
        RECT 38.200 107.900 39.100 108.200 ;
        RECT 34.600 106.900 36.200 107.100 ;
        RECT 35.000 106.800 36.200 106.900 ;
        RECT 37.400 106.800 37.800 107.600 ;
        RECT 31.000 105.800 32.900 106.100 ;
        RECT 24.600 104.800 25.900 105.100 ;
        RECT 24.600 101.100 25.000 104.800 ;
        RECT 25.500 104.700 25.900 104.800 ;
        RECT 26.800 101.100 27.600 105.100 ;
        RECT 28.600 104.800 29.800 105.100 ;
        RECT 28.600 104.700 29.000 104.800 ;
        RECT 29.400 101.100 29.800 104.800 ;
        RECT 31.000 101.100 31.400 105.800 ;
        RECT 32.600 105.200 32.900 105.800 ;
        RECT 31.800 104.400 32.200 105.200 ;
        RECT 32.600 105.100 33.000 105.200 ;
        RECT 33.600 105.100 33.900 106.800 ;
        RECT 34.200 105.800 34.600 106.600 ;
        RECT 32.600 104.800 33.300 105.100 ;
        RECT 33.600 104.800 34.100 105.100 ;
        RECT 33.000 104.200 33.300 104.800 ;
        RECT 33.000 103.800 33.400 104.200 ;
        RECT 33.700 101.100 34.100 104.800 ;
        RECT 35.800 101.100 36.200 106.800 ;
        RECT 37.400 104.100 37.800 104.200 ;
        RECT 38.200 104.100 38.600 107.900 ;
        RECT 41.600 107.100 42.000 109.900 ;
        RECT 46.200 109.200 46.600 109.900 ;
        RECT 46.200 108.800 46.700 109.200 ;
        RECT 47.800 108.900 48.200 109.900 ;
        RECT 47.800 108.800 48.400 108.900 ;
        RECT 46.400 108.500 48.400 108.800 ;
        RECT 43.000 108.100 43.400 108.200 ;
        RECT 44.600 108.100 45.000 108.200 ;
        RECT 45.400 108.100 46.300 108.200 ;
        RECT 43.000 107.800 46.300 108.100 ;
        RECT 43.000 107.100 43.400 107.200 ;
        RECT 46.200 107.100 47.000 107.200 ;
        RECT 41.600 106.900 42.500 107.100 ;
        RECT 41.700 106.800 42.500 106.900 ;
        RECT 43.000 106.800 47.000 107.100 ;
        RECT 40.600 105.800 41.400 106.200 ;
        RECT 39.000 104.400 39.400 105.200 ;
        RECT 39.800 104.800 40.200 105.600 ;
        RECT 42.200 105.200 42.500 106.800 ;
        RECT 47.000 105.800 47.800 106.200 ;
        RECT 48.100 105.200 48.400 108.500 ;
        RECT 51.800 108.200 52.200 109.900 ;
        RECT 51.700 107.900 52.200 108.200 ;
        RECT 51.700 107.200 52.000 107.900 ;
        RECT 53.400 107.600 53.800 109.900 ;
        RECT 52.500 107.300 53.800 107.600 ;
        RECT 54.200 108.500 54.600 109.500 ;
        RECT 54.200 107.400 54.500 108.500 ;
        RECT 56.300 108.000 56.700 109.500 ;
        RECT 60.300 108.200 60.700 109.900 ;
        RECT 56.300 107.700 57.100 108.000 ;
        RECT 56.700 107.500 57.100 107.700 ;
        RECT 59.800 107.900 60.700 108.200 ;
        RECT 61.400 108.000 61.800 109.900 ;
        RECT 63.000 109.600 65.000 109.900 ;
        RECT 63.000 108.000 63.400 109.600 ;
        RECT 61.400 107.900 63.400 108.000 ;
        RECT 63.800 107.900 64.200 109.300 ;
        RECT 64.600 107.900 65.000 109.600 ;
        RECT 66.200 108.900 66.600 109.900 ;
        RECT 51.700 106.800 52.200 107.200 ;
        RECT 42.200 104.800 42.600 105.200 ;
        RECT 48.100 104.900 49.800 105.200 ;
        RECT 49.400 104.800 49.800 104.900 ;
        RECT 51.700 105.100 52.000 106.800 ;
        RECT 52.500 106.500 52.800 107.300 ;
        RECT 54.200 107.100 56.300 107.400 ;
        RECT 55.800 106.900 56.300 107.100 ;
        RECT 56.800 107.200 57.100 107.500 ;
        RECT 52.300 106.100 52.800 106.500 ;
        RECT 52.500 105.100 52.800 106.100 ;
        RECT 53.300 106.200 53.700 106.600 ;
        RECT 53.300 105.800 53.800 106.200 ;
        RECT 54.200 105.800 54.600 106.600 ;
        RECT 55.000 105.800 55.400 106.600 ;
        RECT 55.800 106.500 56.500 106.900 ;
        RECT 56.800 106.800 57.800 107.200 ;
        RECT 59.000 106.800 59.400 107.600 ;
        RECT 55.800 105.500 56.100 106.500 ;
        RECT 54.200 105.200 56.100 105.500 ;
        RECT 37.400 103.800 38.600 104.100 ;
        RECT 41.400 103.800 41.800 104.600 ;
        RECT 38.200 101.100 38.600 103.800 ;
        RECT 42.200 103.500 42.500 104.800 ;
        RECT 44.700 104.400 46.500 104.700 ;
        RECT 44.700 104.100 45.000 104.400 ;
        RECT 40.700 103.200 42.500 103.500 ;
        RECT 40.600 101.100 41.000 103.200 ;
        RECT 42.200 103.100 42.500 103.200 ;
        RECT 42.200 101.100 42.600 103.100 ;
        RECT 44.600 101.100 45.000 104.100 ;
        RECT 46.200 104.100 46.500 104.400 ;
        RECT 47.100 104.500 48.900 104.600 ;
        RECT 49.400 104.500 49.700 104.800 ;
        RECT 51.700 104.600 52.200 105.100 ;
        RECT 52.500 104.800 53.800 105.100 ;
        RECT 47.100 104.300 49.000 104.500 ;
        RECT 47.100 104.100 47.400 104.300 ;
        RECT 46.200 101.400 46.600 104.100 ;
        RECT 47.000 101.700 47.400 104.100 ;
        RECT 47.800 101.400 48.200 104.000 ;
        RECT 48.600 101.500 49.000 104.300 ;
        RECT 49.400 101.700 49.800 104.500 ;
        RECT 46.200 101.100 48.200 101.400 ;
        RECT 48.700 101.400 49.000 101.500 ;
        RECT 50.200 101.500 50.600 104.500 ;
        RECT 50.200 101.400 50.500 101.500 ;
        RECT 48.700 101.100 50.500 101.400 ;
        RECT 51.800 101.100 52.200 104.600 ;
        RECT 53.400 101.100 53.800 104.800 ;
        RECT 54.200 103.500 54.500 105.200 ;
        RECT 56.800 104.900 57.100 106.800 ;
        RECT 57.400 105.400 57.800 106.200 ;
        RECT 56.300 104.600 57.100 104.900 ;
        RECT 59.000 105.100 59.400 105.200 ;
        RECT 59.800 105.100 60.200 107.900 ;
        RECT 61.500 107.700 63.300 107.900 ;
        RECT 61.800 107.200 62.200 107.400 ;
        RECT 63.900 107.200 64.200 107.900 ;
        RECT 65.400 107.800 65.800 108.600 ;
        RECT 66.300 107.200 66.600 108.900 ;
        RECT 67.800 107.900 68.200 109.900 ;
        RECT 69.900 109.200 70.300 109.900 ;
        RECT 69.900 108.800 70.600 109.200 ;
        RECT 69.900 108.400 70.300 108.800 ;
        RECT 69.900 107.900 70.600 108.400 ;
        RECT 71.000 107.900 71.400 109.900 ;
        RECT 71.800 108.000 72.200 109.900 ;
        RECT 73.400 108.000 73.800 109.900 ;
        RECT 71.800 107.900 73.800 108.000 ;
        RECT 67.900 107.800 68.200 107.900 ;
        RECT 67.900 107.600 68.800 107.800 ;
        RECT 67.900 107.500 70.000 107.600 ;
        RECT 68.500 107.300 70.000 107.500 ;
        RECT 69.600 107.200 70.000 107.300 ;
        RECT 61.400 106.900 62.200 107.200 ;
        RECT 63.000 106.900 64.200 107.200 ;
        RECT 61.400 106.800 61.800 106.900 ;
        RECT 63.000 106.800 63.400 106.900 ;
        RECT 62.200 105.800 62.600 106.600 ;
        RECT 59.000 104.800 60.200 105.100 ;
        RECT 54.200 101.500 54.600 103.500 ;
        RECT 56.300 102.200 56.700 104.600 ;
        RECT 55.800 101.800 56.700 102.200 ;
        RECT 56.300 101.100 56.700 101.800 ;
        RECT 59.800 101.100 60.200 104.800 ;
        RECT 60.600 104.400 61.000 105.200 ;
        RECT 63.000 105.100 63.300 106.800 ;
        RECT 63.800 105.800 64.200 106.600 ;
        RECT 64.600 106.400 65.000 107.200 ;
        RECT 66.200 106.800 66.600 107.200 ;
        RECT 65.400 106.100 65.800 106.200 ;
        RECT 66.300 106.100 66.600 106.800 ;
        RECT 67.800 106.400 68.200 107.200 ;
        RECT 68.600 106.600 69.200 107.000 ;
        RECT 68.700 106.200 69.000 106.600 ;
        RECT 65.400 105.800 66.600 106.100 ;
        RECT 66.300 105.100 66.600 105.800 ;
        RECT 67.000 105.400 67.400 106.200 ;
        RECT 68.600 105.800 69.000 106.200 ;
        RECT 69.600 105.500 69.900 107.200 ;
        RECT 70.300 106.200 70.600 107.900 ;
        RECT 71.100 107.200 71.400 107.900 ;
        RECT 71.900 107.700 73.700 107.900 ;
        RECT 73.000 107.200 73.400 107.400 ;
        RECT 71.000 106.800 72.300 107.200 ;
        RECT 73.000 107.100 73.800 107.200 ;
        RECT 74.200 107.100 74.600 109.900 ;
        RECT 75.000 107.800 75.400 108.600 ;
        RECT 76.600 107.600 77.000 109.900 ;
        RECT 78.200 107.600 78.600 109.900 ;
        RECT 79.800 107.600 80.200 109.900 ;
        RECT 81.400 107.600 81.800 109.900 ;
        RECT 73.000 106.900 74.600 107.100 ;
        RECT 73.400 106.800 74.600 106.900 ;
        RECT 70.200 105.800 70.600 106.200 ;
        RECT 68.700 105.200 69.900 105.500 ;
        RECT 62.700 102.200 63.700 105.100 ;
        RECT 66.200 104.700 67.100 105.100 ;
        RECT 62.200 101.800 63.700 102.200 ;
        RECT 62.700 101.100 63.700 101.800 ;
        RECT 66.700 101.100 67.100 104.700 ;
        RECT 68.700 103.100 69.000 105.200 ;
        RECT 70.300 105.100 70.600 105.800 ;
        RECT 68.600 101.100 69.000 103.100 ;
        RECT 70.200 101.100 70.600 105.100 ;
        RECT 71.000 105.100 71.400 105.200 ;
        RECT 72.000 105.100 72.300 106.800 ;
        RECT 72.600 106.100 73.000 106.600 ;
        RECT 73.400 106.100 73.800 106.200 ;
        RECT 72.600 105.800 73.800 106.100 ;
        RECT 71.000 104.800 71.700 105.100 ;
        RECT 72.000 104.800 72.500 105.100 ;
        RECT 71.400 104.200 71.700 104.800 ;
        RECT 71.400 103.800 71.800 104.200 ;
        RECT 72.100 101.100 72.500 104.800 ;
        RECT 74.200 101.100 74.600 106.800 ;
        RECT 75.800 107.200 77.000 107.600 ;
        RECT 77.500 107.200 78.600 107.600 ;
        RECT 79.100 107.200 80.200 107.600 ;
        RECT 80.900 107.200 81.800 107.600 ;
        RECT 83.000 107.700 83.400 109.900 ;
        RECT 85.100 109.200 85.700 109.900 ;
        RECT 85.100 108.900 85.800 109.200 ;
        RECT 87.400 108.900 87.800 109.900 ;
        RECT 89.600 109.200 90.000 109.900 ;
        RECT 89.600 108.900 90.600 109.200 ;
        RECT 85.400 108.500 85.800 108.900 ;
        RECT 87.500 108.600 87.800 108.900 ;
        RECT 87.500 108.300 88.900 108.600 ;
        RECT 88.500 108.200 88.900 108.300 ;
        RECT 89.400 108.200 89.800 108.600 ;
        RECT 90.200 108.500 90.600 108.900 ;
        RECT 84.500 107.700 84.900 107.800 ;
        RECT 83.000 107.400 84.900 107.700 ;
        RECT 75.800 105.800 76.200 107.200 ;
        RECT 77.500 106.900 77.900 107.200 ;
        RECT 79.100 106.900 79.500 107.200 ;
        RECT 80.900 106.900 81.300 107.200 ;
        RECT 76.600 106.500 77.900 106.900 ;
        RECT 78.300 106.500 79.500 106.900 ;
        RECT 80.000 106.500 81.300 106.900 ;
        RECT 77.500 105.800 77.900 106.500 ;
        RECT 79.100 105.800 79.500 106.500 ;
        RECT 80.900 105.800 81.300 106.500 ;
        RECT 75.800 105.400 77.000 105.800 ;
        RECT 77.500 105.400 78.600 105.800 ;
        RECT 79.100 105.400 80.200 105.800 ;
        RECT 80.900 105.400 81.800 105.800 ;
        RECT 76.600 101.100 77.000 105.400 ;
        RECT 78.200 101.100 78.600 105.400 ;
        RECT 79.800 101.100 80.200 105.400 ;
        RECT 81.400 101.100 81.800 105.400 ;
        RECT 83.000 105.700 83.400 107.400 ;
        RECT 86.500 107.100 86.900 107.200 ;
        RECT 89.400 107.100 89.700 108.200 ;
        RECT 91.800 107.500 92.200 109.900 ;
        RECT 94.200 107.700 94.600 109.900 ;
        RECT 96.300 109.200 96.900 109.900 ;
        RECT 96.300 108.900 97.000 109.200 ;
        RECT 98.600 108.900 99.000 109.900 ;
        RECT 100.800 109.200 101.200 109.900 ;
        RECT 100.800 108.900 101.800 109.200 ;
        RECT 96.600 108.500 97.000 108.900 ;
        RECT 98.700 108.600 99.000 108.900 ;
        RECT 98.700 108.300 100.100 108.600 ;
        RECT 99.700 108.200 100.100 108.300 ;
        RECT 100.600 108.200 101.000 108.600 ;
        RECT 101.400 108.500 101.800 108.900 ;
        RECT 95.700 107.700 96.100 107.800 ;
        RECT 94.200 107.400 96.100 107.700 ;
        RECT 91.000 107.100 91.800 107.200 ;
        RECT 86.300 106.800 91.800 107.100 ;
        RECT 85.400 106.400 85.800 106.500 ;
        RECT 83.900 106.100 85.800 106.400 ;
        RECT 83.900 106.000 84.300 106.100 ;
        RECT 84.700 105.700 85.100 105.800 ;
        RECT 83.000 105.400 85.100 105.700 ;
        RECT 83.000 101.100 83.400 105.400 ;
        RECT 86.300 105.200 86.600 106.800 ;
        RECT 89.900 106.700 90.300 106.800 ;
        RECT 89.400 106.200 89.800 106.300 ;
        RECT 90.700 106.200 91.100 106.300 ;
        RECT 88.600 105.900 91.100 106.200 ;
        RECT 88.600 105.800 89.000 105.900 ;
        RECT 94.200 105.700 94.600 107.400 ;
        RECT 97.700 107.100 98.100 107.200 ;
        RECT 99.000 107.100 99.400 107.200 ;
        RECT 100.600 107.100 100.900 108.200 ;
        RECT 103.000 107.500 103.400 109.900 ;
        RECT 103.800 107.700 104.200 109.900 ;
        RECT 105.900 109.200 106.500 109.900 ;
        RECT 105.900 108.900 106.600 109.200 ;
        RECT 108.200 108.900 108.600 109.900 ;
        RECT 110.400 109.200 110.800 109.900 ;
        RECT 110.400 108.900 111.400 109.200 ;
        RECT 106.200 108.500 106.600 108.900 ;
        RECT 108.300 108.600 108.600 108.900 ;
        RECT 108.300 108.300 109.700 108.600 ;
        RECT 109.300 108.200 109.700 108.300 ;
        RECT 110.200 108.200 110.600 108.600 ;
        RECT 111.000 108.500 111.400 108.900 ;
        RECT 105.300 107.700 105.700 107.800 ;
        RECT 103.800 107.400 105.700 107.700 ;
        RECT 102.200 107.100 103.000 107.200 ;
        RECT 97.500 106.800 103.000 107.100 ;
        RECT 96.600 106.400 97.000 106.500 ;
        RECT 95.100 106.100 97.000 106.400 ;
        RECT 95.100 106.000 95.500 106.100 ;
        RECT 95.900 105.700 96.300 105.800 ;
        RECT 89.400 105.500 92.200 105.600 ;
        RECT 89.300 105.400 92.200 105.500 ;
        RECT 85.400 104.900 86.600 105.200 ;
        RECT 87.300 105.300 92.200 105.400 ;
        RECT 87.300 105.100 89.700 105.300 ;
        RECT 85.400 104.400 85.700 104.900 ;
        RECT 85.000 104.000 85.700 104.400 ;
        RECT 86.500 104.500 86.900 104.600 ;
        RECT 87.300 104.500 87.600 105.100 ;
        RECT 86.500 104.200 87.600 104.500 ;
        RECT 87.900 104.500 90.600 104.800 ;
        RECT 87.900 104.400 88.300 104.500 ;
        RECT 90.200 104.400 90.600 104.500 ;
        RECT 87.100 103.700 87.500 103.800 ;
        RECT 88.500 103.700 88.900 103.800 ;
        RECT 85.400 103.100 85.800 103.500 ;
        RECT 87.100 103.400 88.900 103.700 ;
        RECT 87.500 103.100 87.800 103.400 ;
        RECT 90.200 103.100 90.600 103.500 ;
        RECT 85.100 101.100 85.700 103.100 ;
        RECT 87.400 101.100 87.800 103.100 ;
        RECT 89.600 102.800 90.600 103.100 ;
        RECT 89.600 101.100 90.000 102.800 ;
        RECT 91.800 101.100 92.200 105.300 ;
        RECT 94.200 105.400 96.300 105.700 ;
        RECT 94.200 101.100 94.600 105.400 ;
        RECT 97.500 105.200 97.800 106.800 ;
        RECT 101.100 106.700 101.500 106.800 ;
        RECT 101.900 106.200 102.300 106.300 ;
        RECT 99.800 105.900 102.300 106.200 ;
        RECT 99.800 105.800 100.200 105.900 ;
        RECT 103.800 105.700 104.200 107.400 ;
        RECT 107.300 107.100 107.700 107.200 ;
        RECT 110.200 107.100 110.500 108.200 ;
        RECT 112.600 107.500 113.000 109.900 ;
        RECT 114.200 108.900 114.600 109.900 ;
        RECT 113.400 107.800 113.800 108.600 ;
        RECT 114.300 107.200 114.600 108.900 ;
        RECT 116.600 107.600 117.000 109.900 ;
        RECT 118.200 107.600 118.600 109.900 ;
        RECT 119.800 107.600 120.200 109.900 ;
        RECT 121.400 107.600 121.800 109.900 ;
        RECT 111.800 107.100 112.600 107.200 ;
        RECT 107.100 106.800 112.600 107.100 ;
        RECT 113.400 106.800 113.800 107.200 ;
        RECT 114.200 106.800 114.600 107.200 ;
        RECT 106.200 106.400 106.600 106.500 ;
        RECT 104.700 106.100 106.600 106.400 ;
        RECT 107.100 106.200 107.400 106.800 ;
        RECT 110.700 106.700 111.100 106.800 ;
        RECT 110.200 106.200 110.600 106.300 ;
        RECT 111.500 106.200 111.900 106.300 ;
        RECT 104.700 106.000 105.100 106.100 ;
        RECT 107.000 105.800 107.400 106.200 ;
        RECT 109.400 105.900 111.900 106.200 ;
        RECT 113.400 106.100 113.700 106.800 ;
        RECT 114.300 106.100 114.600 106.800 ;
        RECT 115.800 107.200 117.000 107.600 ;
        RECT 117.500 107.200 118.600 107.600 ;
        RECT 119.100 107.200 120.200 107.600 ;
        RECT 120.900 107.200 121.800 107.600 ;
        RECT 123.000 108.500 123.400 109.500 ;
        RECT 123.000 107.400 123.300 108.500 ;
        RECT 125.100 108.000 125.500 109.500 ;
        RECT 125.100 107.700 125.900 108.000 ;
        RECT 125.500 107.500 125.900 107.700 ;
        RECT 127.800 107.500 128.200 109.900 ;
        RECT 130.000 109.200 130.400 109.900 ;
        RECT 129.400 108.900 130.400 109.200 ;
        RECT 132.200 108.900 132.600 109.900 ;
        RECT 134.300 109.200 134.900 109.900 ;
        RECT 134.200 108.900 134.900 109.200 ;
        RECT 129.400 108.500 129.800 108.900 ;
        RECT 132.200 108.600 132.500 108.900 ;
        RECT 130.200 108.200 130.600 108.600 ;
        RECT 131.100 108.300 132.500 108.600 ;
        RECT 134.200 108.500 134.600 108.900 ;
        RECT 131.100 108.200 131.500 108.300 ;
        RECT 109.400 105.800 109.800 105.900 ;
        RECT 113.400 105.800 114.600 106.100 ;
        RECT 105.500 105.700 105.900 105.800 ;
        RECT 100.600 105.500 103.400 105.600 ;
        RECT 100.500 105.400 103.400 105.500 ;
        RECT 96.600 104.900 97.800 105.200 ;
        RECT 98.500 105.300 103.400 105.400 ;
        RECT 98.500 105.100 100.900 105.300 ;
        RECT 96.600 104.400 96.900 104.900 ;
        RECT 96.200 104.000 96.900 104.400 ;
        RECT 97.700 104.500 98.100 104.600 ;
        RECT 98.500 104.500 98.800 105.100 ;
        RECT 97.700 104.200 98.800 104.500 ;
        RECT 99.100 104.500 101.800 104.800 ;
        RECT 99.100 104.400 99.500 104.500 ;
        RECT 101.400 104.400 101.800 104.500 ;
        RECT 98.300 103.700 98.700 103.800 ;
        RECT 99.700 103.700 100.100 103.800 ;
        RECT 96.600 103.100 97.000 103.500 ;
        RECT 98.300 103.400 100.100 103.700 ;
        RECT 98.700 103.100 99.000 103.400 ;
        RECT 101.400 103.100 101.800 103.500 ;
        RECT 96.300 101.100 96.900 103.100 ;
        RECT 98.600 101.100 99.000 103.100 ;
        RECT 100.800 102.800 101.800 103.100 ;
        RECT 100.800 101.100 101.200 102.800 ;
        RECT 103.000 101.100 103.400 105.300 ;
        RECT 103.800 105.400 105.900 105.700 ;
        RECT 103.800 101.100 104.200 105.400 ;
        RECT 107.100 105.200 107.400 105.800 ;
        RECT 110.200 105.500 113.000 105.600 ;
        RECT 110.100 105.400 113.000 105.500 ;
        RECT 106.200 104.900 107.400 105.200 ;
        RECT 108.100 105.300 113.000 105.400 ;
        RECT 108.100 105.100 110.500 105.300 ;
        RECT 106.200 104.400 106.500 104.900 ;
        RECT 105.800 104.000 106.500 104.400 ;
        RECT 107.300 104.500 107.700 104.600 ;
        RECT 108.100 104.500 108.400 105.100 ;
        RECT 107.300 104.200 108.400 104.500 ;
        RECT 108.700 104.500 111.400 104.800 ;
        RECT 108.700 104.400 109.100 104.500 ;
        RECT 111.000 104.400 111.400 104.500 ;
        RECT 107.900 103.700 108.300 103.800 ;
        RECT 109.300 103.700 109.700 103.800 ;
        RECT 106.200 103.100 106.600 103.500 ;
        RECT 107.900 103.400 109.700 103.700 ;
        RECT 108.300 103.100 108.600 103.400 ;
        RECT 111.000 103.100 111.400 103.500 ;
        RECT 105.900 101.100 106.500 103.100 ;
        RECT 108.200 101.100 108.600 103.100 ;
        RECT 110.400 102.800 111.400 103.100 ;
        RECT 110.400 101.100 110.800 102.800 ;
        RECT 112.600 101.100 113.000 105.300 ;
        RECT 114.300 105.100 114.600 105.800 ;
        RECT 115.000 105.400 115.400 106.200 ;
        RECT 115.800 105.800 116.200 107.200 ;
        RECT 117.500 106.900 117.900 107.200 ;
        RECT 119.100 106.900 119.500 107.200 ;
        RECT 120.900 106.900 121.300 107.200 ;
        RECT 123.000 107.100 125.100 107.400 ;
        RECT 116.600 106.500 117.900 106.900 ;
        RECT 118.300 106.500 119.500 106.900 ;
        RECT 120.000 106.500 121.300 106.900 ;
        RECT 124.600 106.900 125.100 107.100 ;
        RECT 125.600 107.200 125.900 107.500 ;
        RECT 117.500 105.800 117.900 106.500 ;
        RECT 119.100 105.800 119.500 106.500 ;
        RECT 120.900 105.800 121.300 106.500 ;
        RECT 123.000 105.800 123.400 106.600 ;
        RECT 123.800 105.800 124.200 106.600 ;
        RECT 124.600 106.500 125.300 106.900 ;
        RECT 125.600 106.800 126.600 107.200 ;
        RECT 128.200 107.100 129.000 107.200 ;
        RECT 130.300 107.100 130.600 108.200 ;
        RECT 135.100 107.700 135.500 107.800 ;
        RECT 136.600 107.700 137.000 109.900 ;
        RECT 135.100 107.400 137.000 107.700 ;
        RECT 137.400 107.500 137.800 109.900 ;
        RECT 139.600 109.200 140.000 109.900 ;
        RECT 139.000 108.900 140.000 109.200 ;
        RECT 141.800 108.900 142.200 109.900 ;
        RECT 143.900 109.200 144.500 109.900 ;
        RECT 143.800 108.900 144.500 109.200 ;
        RECT 139.000 108.500 139.400 108.900 ;
        RECT 141.800 108.600 142.100 108.900 ;
        RECT 139.800 108.200 140.200 108.600 ;
        RECT 140.700 108.300 142.100 108.600 ;
        RECT 143.800 108.500 144.200 108.900 ;
        RECT 140.700 108.200 141.100 108.300 ;
        RECT 133.100 107.100 133.500 107.200 ;
        RECT 128.200 106.800 133.700 107.100 ;
        RECT 115.800 105.400 117.000 105.800 ;
        RECT 117.500 105.400 118.600 105.800 ;
        RECT 119.100 105.400 120.200 105.800 ;
        RECT 120.900 105.400 121.800 105.800 ;
        RECT 124.600 105.500 124.900 106.500 ;
        RECT 114.200 104.700 115.100 105.100 ;
        RECT 114.700 101.100 115.100 104.700 ;
        RECT 116.600 101.100 117.000 105.400 ;
        RECT 118.200 101.100 118.600 105.400 ;
        RECT 119.800 101.100 120.200 105.400 ;
        RECT 121.400 101.100 121.800 105.400 ;
        RECT 123.000 105.200 124.900 105.500 ;
        RECT 123.000 103.500 123.300 105.200 ;
        RECT 125.600 104.900 125.900 106.800 ;
        RECT 129.700 106.700 130.100 106.800 ;
        RECT 128.900 106.200 129.300 106.300 ;
        RECT 126.200 105.400 126.600 106.200 ;
        RECT 128.900 105.900 131.400 106.200 ;
        RECT 131.000 105.800 131.400 105.900 ;
        RECT 127.800 105.500 130.600 105.600 ;
        RECT 127.800 105.400 130.700 105.500 ;
        RECT 125.100 104.600 125.900 104.900 ;
        RECT 127.800 105.300 132.700 105.400 ;
        RECT 123.000 101.500 123.400 103.500 ;
        RECT 125.100 102.200 125.500 104.600 ;
        RECT 125.100 101.800 125.800 102.200 ;
        RECT 125.100 101.100 125.500 101.800 ;
        RECT 127.800 101.100 128.200 105.300 ;
        RECT 130.300 105.100 132.700 105.300 ;
        RECT 129.400 104.500 132.100 104.800 ;
        RECT 129.400 104.400 129.800 104.500 ;
        RECT 131.700 104.400 132.100 104.500 ;
        RECT 132.400 104.500 132.700 105.100 ;
        RECT 133.400 105.200 133.700 106.800 ;
        RECT 134.200 106.400 134.600 106.500 ;
        RECT 134.200 106.100 136.100 106.400 ;
        RECT 135.700 106.000 136.100 106.100 ;
        RECT 134.900 105.700 135.300 105.800 ;
        RECT 136.600 105.700 137.000 107.400 ;
        RECT 137.800 107.100 138.600 107.200 ;
        RECT 139.900 107.100 140.200 108.200 ;
        RECT 144.700 107.700 145.100 107.800 ;
        RECT 146.200 107.700 146.600 109.900 ;
        RECT 148.300 108.200 148.700 109.900 ;
        RECT 144.700 107.400 146.600 107.700 ;
        RECT 147.800 107.900 148.700 108.200 ;
        RECT 151.000 107.900 151.400 109.900 ;
        RECT 151.800 108.000 152.200 109.900 ;
        RECT 153.400 108.000 153.800 109.900 ;
        RECT 151.800 107.900 153.800 108.000 ;
        RECT 142.700 107.100 143.100 107.200 ;
        RECT 137.800 106.800 143.300 107.100 ;
        RECT 139.300 106.700 139.700 106.800 ;
        RECT 138.500 106.200 138.900 106.300 ;
        RECT 138.500 106.100 141.000 106.200 ;
        RECT 141.400 106.100 141.800 106.200 ;
        RECT 138.500 105.900 141.800 106.100 ;
        RECT 140.600 105.800 141.800 105.900 ;
        RECT 134.900 105.400 137.000 105.700 ;
        RECT 133.400 104.900 134.600 105.200 ;
        RECT 133.100 104.500 133.500 104.600 ;
        RECT 132.400 104.200 133.500 104.500 ;
        RECT 134.300 104.400 134.600 104.900 ;
        RECT 134.300 104.000 135.000 104.400 ;
        RECT 131.100 103.700 131.500 103.800 ;
        RECT 132.500 103.700 132.900 103.800 ;
        RECT 129.400 103.100 129.800 103.500 ;
        RECT 131.100 103.400 132.900 103.700 ;
        RECT 132.200 103.100 132.500 103.400 ;
        RECT 134.200 103.100 134.600 103.500 ;
        RECT 129.400 102.800 130.400 103.100 ;
        RECT 130.000 101.100 130.400 102.800 ;
        RECT 132.200 101.100 132.600 103.100 ;
        RECT 134.300 101.100 134.900 103.100 ;
        RECT 136.600 101.100 137.000 105.400 ;
        RECT 137.400 105.500 140.200 105.600 ;
        RECT 137.400 105.400 140.300 105.500 ;
        RECT 137.400 105.300 142.300 105.400 ;
        RECT 137.400 101.100 137.800 105.300 ;
        RECT 139.900 105.100 142.300 105.300 ;
        RECT 139.000 104.500 141.700 104.800 ;
        RECT 139.000 104.400 139.400 104.500 ;
        RECT 141.300 104.400 141.700 104.500 ;
        RECT 142.000 104.500 142.300 105.100 ;
        RECT 143.000 105.200 143.300 106.800 ;
        RECT 143.800 106.400 144.200 106.500 ;
        RECT 143.800 106.100 145.700 106.400 ;
        RECT 145.300 106.000 145.700 106.100 ;
        RECT 144.500 105.700 144.900 105.800 ;
        RECT 146.200 105.700 146.600 107.400 ;
        RECT 147.000 106.800 147.400 107.600 ;
        RECT 144.500 105.400 146.600 105.700 ;
        RECT 143.000 104.900 144.200 105.200 ;
        RECT 142.700 104.500 143.100 104.600 ;
        RECT 142.000 104.200 143.100 104.500 ;
        RECT 143.900 104.400 144.200 104.900 ;
        RECT 143.900 104.000 144.600 104.400 ;
        RECT 140.700 103.700 141.100 103.800 ;
        RECT 142.100 103.700 142.500 103.800 ;
        RECT 139.000 103.100 139.400 103.500 ;
        RECT 140.700 103.400 142.500 103.700 ;
        RECT 141.800 103.100 142.100 103.400 ;
        RECT 143.800 103.100 144.200 103.500 ;
        RECT 139.000 102.800 140.000 103.100 ;
        RECT 139.600 101.100 140.000 102.800 ;
        RECT 141.800 101.100 142.200 103.100 ;
        RECT 143.900 101.100 144.500 103.100 ;
        RECT 146.200 101.100 146.600 105.400 ;
        RECT 147.800 106.100 148.200 107.900 ;
        RECT 151.100 107.200 151.400 107.900 ;
        RECT 151.900 107.700 153.700 107.900 ;
        RECT 153.000 107.200 153.400 107.400 ;
        RECT 151.000 106.800 152.300 107.200 ;
        RECT 153.000 107.100 153.800 107.200 ;
        RECT 154.200 107.100 154.600 109.900 ;
        RECT 156.600 108.900 157.000 109.900 ;
        RECT 155.000 107.800 155.400 108.600 ;
        RECT 155.800 107.800 156.200 108.600 ;
        RECT 156.700 107.200 157.000 108.900 ;
        RECT 158.200 109.600 160.200 109.900 ;
        RECT 158.200 107.900 158.600 109.600 ;
        RECT 159.000 107.900 159.400 109.300 ;
        RECT 159.800 108.000 160.200 109.600 ;
        RECT 161.400 108.000 161.800 109.900 ;
        RECT 163.000 108.900 163.400 109.900 ;
        RECT 164.900 109.200 165.300 109.900 ;
        RECT 159.800 107.900 161.800 108.000 ;
        RECT 159.000 107.200 159.300 107.900 ;
        RECT 159.900 107.700 161.700 107.900 ;
        RECT 162.200 107.800 162.600 108.600 ;
        RECT 161.000 107.200 161.400 107.400 ;
        RECT 163.100 107.200 163.400 108.900 ;
        RECT 164.600 108.800 165.300 109.200 ;
        RECT 164.900 108.400 165.300 108.800 ;
        RECT 153.000 106.900 154.600 107.100 ;
        RECT 153.400 106.800 154.600 106.900 ;
        RECT 156.600 106.800 157.000 107.200 ;
        RECT 147.800 105.800 151.300 106.100 ;
        RECT 147.800 101.100 148.200 105.800 ;
        RECT 151.000 105.200 151.300 105.800 ;
        RECT 148.600 105.100 149.000 105.200 ;
        RECT 149.400 105.100 149.800 105.200 ;
        RECT 148.600 104.800 149.800 105.100 ;
        RECT 151.000 105.100 151.400 105.200 ;
        RECT 152.000 105.100 152.300 106.800 ;
        RECT 152.600 105.800 153.000 106.600 ;
        RECT 151.000 104.800 151.700 105.100 ;
        RECT 152.000 104.800 152.500 105.100 ;
        RECT 148.600 104.400 149.000 104.800 ;
        RECT 151.400 104.200 151.700 104.800 ;
        RECT 151.400 103.800 151.800 104.200 ;
        RECT 152.100 101.100 152.500 104.800 ;
        RECT 154.200 101.100 154.600 106.800 ;
        RECT 155.800 106.100 156.200 106.200 ;
        RECT 156.700 106.100 157.000 106.800 ;
        RECT 158.200 106.400 158.600 107.200 ;
        RECT 159.000 106.900 160.200 107.200 ;
        RECT 161.000 106.900 161.800 107.200 ;
        RECT 159.800 106.800 160.200 106.900 ;
        RECT 161.400 106.800 161.800 106.900 ;
        RECT 163.000 106.800 163.400 107.200 ;
        RECT 155.800 105.800 157.000 106.100 ;
        RECT 156.700 105.100 157.000 105.800 ;
        RECT 157.400 105.400 157.800 106.200 ;
        RECT 159.000 105.800 159.400 106.600 ;
        RECT 159.900 105.100 160.200 106.800 ;
        RECT 160.600 106.100 161.000 106.600 ;
        RECT 163.100 106.100 163.400 106.800 ;
        RECT 164.600 107.900 165.300 108.400 ;
        RECT 167.000 107.900 167.400 109.900 ;
        RECT 167.800 108.500 168.200 109.500 ;
        RECT 164.600 106.200 164.900 107.900 ;
        RECT 167.000 107.800 167.300 107.900 ;
        RECT 166.400 107.600 167.300 107.800 ;
        RECT 165.200 107.500 167.300 107.600 ;
        RECT 165.200 107.300 166.700 107.500 ;
        RECT 167.800 107.400 168.100 108.500 ;
        RECT 169.900 108.000 170.300 109.500 ;
        RECT 173.400 108.800 173.800 109.900 ;
        RECT 169.900 107.700 170.700 108.000 ;
        RECT 170.300 107.500 170.700 107.700 ;
        RECT 165.200 107.200 165.600 107.300 ;
        RECT 160.600 105.800 163.400 106.100 ;
        RECT 163.100 105.100 163.400 105.800 ;
        RECT 163.800 105.400 164.200 106.200 ;
        RECT 164.600 105.800 165.000 106.200 ;
        RECT 164.600 105.100 164.900 105.800 ;
        RECT 165.300 105.500 165.600 107.200 ;
        RECT 166.000 106.900 166.400 107.000 ;
        RECT 166.000 106.600 166.500 106.900 ;
        RECT 166.200 106.200 166.500 106.600 ;
        RECT 167.000 106.400 167.400 107.200 ;
        RECT 167.800 107.100 169.900 107.400 ;
        RECT 169.400 106.900 169.900 107.100 ;
        RECT 170.400 107.200 170.700 107.500 ;
        RECT 173.400 107.200 173.700 108.800 ;
        RECT 174.200 107.800 174.600 108.600 ;
        RECT 175.800 107.600 176.200 109.900 ;
        RECT 177.400 107.600 177.800 109.900 ;
        RECT 179.000 107.600 179.400 109.900 ;
        RECT 180.600 107.600 181.000 109.900 ;
        RECT 184.100 109.200 184.500 109.500 ;
        RECT 184.100 108.800 185.000 109.200 ;
        RECT 184.100 108.000 184.500 108.800 ;
        RECT 186.200 108.500 186.600 109.500 ;
        RECT 183.700 107.700 184.500 108.000 ;
        RECT 175.800 107.200 176.700 107.600 ;
        RECT 177.400 107.200 178.500 107.600 ;
        RECT 179.000 107.200 180.100 107.600 ;
        RECT 180.600 107.200 181.800 107.600 ;
        RECT 183.700 107.500 184.100 107.700 ;
        RECT 183.700 107.200 184.000 107.500 ;
        RECT 186.300 107.400 186.600 108.500 ;
        RECT 170.400 107.100 171.400 107.200 ;
        RECT 166.200 105.800 166.600 106.200 ;
        RECT 167.800 105.800 168.200 106.600 ;
        RECT 168.600 105.800 169.000 106.600 ;
        RECT 169.400 106.500 170.100 106.900 ;
        RECT 170.400 106.800 172.900 107.100 ;
        RECT 169.400 105.500 169.700 106.500 ;
        RECT 165.300 105.200 166.500 105.500 ;
        RECT 156.600 104.700 157.500 105.100 ;
        RECT 157.100 101.100 157.500 104.700 ;
        RECT 159.500 102.200 160.500 105.100 ;
        RECT 163.000 104.700 163.900 105.100 ;
        RECT 159.000 101.800 160.500 102.200 ;
        RECT 159.500 101.100 160.500 101.800 ;
        RECT 163.500 101.100 163.900 104.700 ;
        RECT 164.600 101.100 165.000 105.100 ;
        RECT 166.200 103.100 166.500 105.200 ;
        RECT 167.800 105.200 169.700 105.500 ;
        RECT 167.800 103.500 168.100 105.200 ;
        RECT 170.400 104.900 170.700 106.800 ;
        RECT 172.600 106.200 172.900 106.800 ;
        RECT 173.400 106.800 173.800 107.200 ;
        RECT 176.300 106.900 176.700 107.200 ;
        RECT 178.100 106.900 178.500 107.200 ;
        RECT 179.700 106.900 180.100 107.200 ;
        RECT 171.000 106.100 171.400 106.200 ;
        RECT 171.800 106.100 172.200 106.200 ;
        RECT 171.000 105.800 172.200 106.100 ;
        RECT 171.000 105.400 171.400 105.800 ;
        RECT 172.600 105.400 173.000 106.200 ;
        RECT 173.400 105.100 173.700 106.800 ;
        RECT 176.300 106.500 177.600 106.900 ;
        RECT 178.100 106.500 179.300 106.900 ;
        RECT 179.700 106.500 181.000 106.900 ;
        RECT 176.300 105.800 176.700 106.500 ;
        RECT 178.100 105.800 178.500 106.500 ;
        RECT 179.700 105.800 180.100 106.500 ;
        RECT 181.400 105.800 181.800 107.200 ;
        RECT 183.000 106.800 184.000 107.200 ;
        RECT 184.500 107.100 186.600 107.400 ;
        RECT 187.000 108.500 187.400 109.500 ;
        RECT 189.100 109.200 189.500 109.500 ;
        RECT 189.100 108.800 189.800 109.200 ;
        RECT 192.600 108.900 193.000 109.900 ;
        RECT 187.000 107.400 187.300 108.500 ;
        RECT 189.100 108.000 189.500 108.800 ;
        RECT 189.100 107.700 189.900 108.000 ;
        RECT 191.800 107.800 192.200 108.600 ;
        RECT 192.700 107.800 193.000 108.900 ;
        RECT 194.200 107.900 194.600 109.900 ;
        RECT 189.500 107.500 189.900 107.700 ;
        RECT 192.700 107.500 193.900 107.800 ;
        RECT 187.000 107.100 189.100 107.400 ;
        RECT 184.500 106.900 185.000 107.100 ;
        RECT 175.800 105.400 176.700 105.800 ;
        RECT 177.400 105.400 178.500 105.800 ;
        RECT 179.000 105.400 180.100 105.800 ;
        RECT 180.600 105.400 181.800 105.800 ;
        RECT 183.000 105.400 183.400 106.200 ;
        RECT 169.900 104.600 170.700 104.900 ;
        RECT 172.900 104.700 173.800 105.100 ;
        RECT 166.200 101.100 166.600 103.100 ;
        RECT 167.800 101.500 168.200 103.500 ;
        RECT 169.900 101.100 170.300 104.600 ;
        RECT 172.900 101.100 173.300 104.700 ;
        RECT 175.800 101.100 176.200 105.400 ;
        RECT 177.400 101.100 177.800 105.400 ;
        RECT 179.000 101.100 179.400 105.400 ;
        RECT 180.600 101.100 181.000 105.400 ;
        RECT 183.700 104.900 184.000 106.800 ;
        RECT 184.300 106.500 185.000 106.900 ;
        RECT 188.600 106.900 189.100 107.100 ;
        RECT 189.600 107.200 189.900 107.500 ;
        RECT 184.700 105.500 185.000 106.500 ;
        RECT 185.400 105.800 185.800 106.600 ;
        RECT 186.200 106.100 186.600 106.600 ;
        RECT 187.000 106.100 187.400 106.600 ;
        RECT 186.200 105.800 187.400 106.100 ;
        RECT 187.800 105.800 188.200 106.600 ;
        RECT 188.600 106.500 189.300 106.900 ;
        RECT 189.600 106.800 190.600 107.200 ;
        RECT 192.600 106.800 193.100 107.200 ;
        RECT 188.600 105.500 188.900 106.500 ;
        RECT 184.700 105.200 186.600 105.500 ;
        RECT 183.700 104.600 184.500 104.900 ;
        RECT 184.100 101.100 184.500 104.600 ;
        RECT 186.300 103.500 186.600 105.200 ;
        RECT 186.200 101.500 186.600 103.500 ;
        RECT 187.000 105.200 188.900 105.500 ;
        RECT 187.000 103.500 187.300 105.200 ;
        RECT 189.600 104.900 189.900 106.800 ;
        RECT 192.800 106.400 193.200 106.800 ;
        RECT 190.200 105.400 190.600 106.200 ;
        RECT 193.600 106.000 193.900 107.500 ;
        RECT 194.300 106.200 194.600 107.900 ;
        RECT 193.500 105.700 193.900 106.000 ;
        RECT 194.200 105.800 194.600 106.200 ;
        RECT 191.800 105.600 193.900 105.700 ;
        RECT 191.800 105.400 193.800 105.600 ;
        RECT 189.100 104.600 189.900 104.900 ;
        RECT 187.000 101.500 187.400 103.500 ;
        RECT 189.100 101.100 189.500 104.600 ;
        RECT 191.800 101.100 192.200 105.400 ;
        RECT 194.300 105.100 194.600 105.800 ;
        RECT 193.900 104.800 194.600 105.100 ;
        RECT 193.900 101.100 194.300 104.800 ;
        RECT 2.200 96.200 2.600 99.900 ;
        RECT 3.400 96.800 3.800 97.200 ;
        RECT 3.400 96.200 3.700 96.800 ;
        RECT 4.100 96.200 4.500 99.900 ;
        RECT 1.500 95.900 2.600 96.200 ;
        RECT 3.000 95.900 3.700 96.200 ;
        RECT 4.000 95.900 4.500 96.200 ;
        RECT 1.500 95.600 1.800 95.900 ;
        RECT 3.000 95.800 3.400 95.900 ;
        RECT 1.200 95.200 1.800 95.600 ;
        RECT 1.500 93.700 1.800 95.200 ;
        RECT 2.200 95.100 2.600 95.200 ;
        RECT 3.000 95.100 3.400 95.200 ;
        RECT 2.200 94.800 3.400 95.100 ;
        RECT 2.200 94.400 2.600 94.800 ;
        RECT 4.000 94.200 4.300 95.900 ;
        RECT 4.600 95.100 5.000 95.200 ;
        RECT 5.400 95.100 5.800 95.200 ;
        RECT 4.600 94.800 5.800 95.100 ;
        RECT 4.600 94.400 5.000 94.800 ;
        RECT 3.000 93.800 4.300 94.200 ;
        RECT 5.400 94.100 5.800 94.200 ;
        RECT 6.200 94.100 6.600 99.900 ;
        RECT 7.800 96.200 8.200 99.900 ;
        RECT 8.700 96.200 9.100 96.300 ;
        RECT 7.800 95.900 9.100 96.200 ;
        RECT 10.000 95.900 10.800 99.900 ;
        RECT 11.800 96.200 12.200 96.300 ;
        RECT 12.600 96.200 13.000 99.900 ;
        RECT 11.800 95.900 13.000 96.200 ;
        RECT 9.300 95.200 9.700 95.300 ;
        RECT 10.300 95.200 10.600 95.900 ;
        RECT 8.900 94.900 9.700 95.200 ;
        RECT 8.900 94.800 9.300 94.900 ;
        RECT 10.200 94.800 10.600 95.200 ;
        RECT 9.600 94.300 10.000 94.400 ;
        RECT 8.600 94.200 10.000 94.300 ;
        RECT 5.000 93.800 6.600 94.100 ;
        RECT 7.000 94.100 7.400 94.200 ;
        RECT 7.800 94.100 10.000 94.200 ;
        RECT 7.000 94.000 10.000 94.100 ;
        RECT 10.300 94.200 10.600 94.800 ;
        RECT 13.400 95.600 13.800 99.900 ;
        RECT 15.500 97.900 16.100 99.900 ;
        RECT 17.800 97.900 18.200 99.900 ;
        RECT 20.000 98.200 20.400 99.900 ;
        RECT 20.000 97.900 21.000 98.200 ;
        RECT 15.800 97.500 16.200 97.900 ;
        RECT 17.900 97.600 18.200 97.900 ;
        RECT 17.500 97.300 19.300 97.600 ;
        RECT 20.600 97.500 21.000 97.900 ;
        RECT 17.500 97.200 17.900 97.300 ;
        RECT 18.900 97.200 19.300 97.300 ;
        RECT 15.400 96.600 16.100 97.000 ;
        RECT 15.800 96.100 16.100 96.600 ;
        RECT 16.900 96.500 18.000 96.800 ;
        RECT 16.900 96.400 17.300 96.500 ;
        RECT 15.800 95.800 17.000 96.100 ;
        RECT 13.400 95.300 15.500 95.600 ;
        RECT 7.000 93.900 8.900 94.000 ;
        RECT 10.300 93.900 10.800 94.200 ;
        RECT 7.000 93.800 8.600 93.900 ;
        RECT 1.500 93.400 2.600 93.700 ;
        RECT 2.200 91.100 2.600 93.400 ;
        RECT 3.100 93.100 3.400 93.800 ;
        RECT 5.000 93.600 5.400 93.800 ;
        RECT 3.900 93.100 5.700 93.300 ;
        RECT 3.000 91.100 3.400 93.100 ;
        RECT 3.800 93.000 5.800 93.100 ;
        RECT 3.800 91.100 4.200 93.000 ;
        RECT 5.400 91.100 5.800 93.000 ;
        RECT 6.200 91.100 6.600 93.800 ;
        RECT 8.700 93.400 9.100 93.500 ;
        RECT 7.000 92.400 7.400 93.200 ;
        RECT 7.800 93.100 9.100 93.400 ;
        RECT 9.400 93.200 10.200 93.600 ;
        RECT 7.800 91.100 8.200 93.100 ;
        RECT 10.500 92.900 10.800 93.900 ;
        RECT 11.200 93.800 11.600 94.200 ;
        RECT 12.200 94.100 13.000 94.200 ;
        RECT 13.400 94.100 13.800 95.300 ;
        RECT 15.100 95.200 15.500 95.300 ;
        RECT 16.700 95.200 17.000 95.800 ;
        RECT 17.700 95.900 18.000 96.500 ;
        RECT 18.300 96.500 18.700 96.600 ;
        RECT 20.600 96.500 21.000 96.600 ;
        RECT 18.300 96.200 21.000 96.500 ;
        RECT 17.700 95.700 20.100 95.900 ;
        RECT 22.200 95.700 22.600 99.900 ;
        RECT 23.100 99.600 24.900 99.900 ;
        RECT 23.100 99.500 23.400 99.600 ;
        RECT 23.000 96.500 23.400 99.500 ;
        RECT 24.600 99.500 24.900 99.600 ;
        RECT 25.400 99.600 27.400 99.900 ;
        RECT 23.800 96.500 24.200 99.300 ;
        RECT 24.600 96.700 25.000 99.500 ;
        RECT 25.400 97.000 25.800 99.600 ;
        RECT 26.200 96.900 26.600 99.300 ;
        RECT 27.000 96.900 27.400 99.600 ;
        RECT 26.200 96.700 26.500 96.900 ;
        RECT 24.600 96.500 26.500 96.700 ;
        RECT 23.900 96.200 24.200 96.500 ;
        RECT 24.700 96.400 26.500 96.500 ;
        RECT 27.100 96.600 27.400 96.900 ;
        RECT 28.600 96.900 29.000 99.900 ;
        RECT 28.600 96.600 28.900 96.900 ;
        RECT 27.100 96.300 28.900 96.600 ;
        RECT 23.800 96.100 24.200 96.200 ;
        RECT 23.800 95.800 25.500 96.100 ;
        RECT 29.400 95.900 29.800 99.900 ;
        RECT 30.200 96.200 30.600 99.900 ;
        RECT 31.800 96.200 32.200 99.900 ;
        RECT 30.200 95.900 32.200 96.200 ;
        RECT 33.900 96.200 34.300 99.900 ;
        RECT 34.600 96.800 35.000 97.200 ;
        RECT 34.700 96.200 35.000 96.800 ;
        RECT 37.100 96.200 37.500 99.900 ;
        RECT 37.800 96.800 38.200 97.200 ;
        RECT 37.900 96.200 38.200 96.800 ;
        RECT 39.300 96.300 39.700 99.900 ;
        RECT 33.900 95.900 34.400 96.200 ;
        RECT 34.700 95.900 35.400 96.200 ;
        RECT 37.100 95.900 37.600 96.200 ;
        RECT 37.900 95.900 38.600 96.200 ;
        RECT 39.300 95.900 40.200 96.300 ;
        RECT 17.700 95.600 22.600 95.700 ;
        RECT 19.700 95.500 22.600 95.600 ;
        RECT 19.800 95.400 22.600 95.500 ;
        RECT 14.300 94.900 14.700 95.000 ;
        RECT 14.300 94.600 16.200 94.900 ;
        RECT 16.600 94.800 17.000 95.200 ;
        RECT 19.000 95.100 19.400 95.200 ;
        RECT 19.000 94.800 21.500 95.100 ;
        RECT 15.800 94.500 16.200 94.600 ;
        RECT 12.200 93.800 13.800 94.100 ;
        RECT 16.700 94.200 17.000 94.800 ;
        RECT 19.800 94.700 20.200 94.800 ;
        RECT 21.100 94.700 21.500 94.800 ;
        RECT 20.300 94.200 20.700 94.300 ;
        RECT 25.200 94.200 25.500 95.800 ;
        RECT 29.500 95.200 29.800 95.900 ;
        RECT 31.400 95.200 31.800 95.400 ;
        RECT 25.800 94.800 26.600 95.200 ;
        RECT 28.600 95.100 29.000 95.200 ;
        RECT 29.400 95.100 30.600 95.200 ;
        RECT 28.600 94.900 30.600 95.100 ;
        RECT 31.400 95.100 32.200 95.200 ;
        RECT 31.400 94.900 32.900 95.100 ;
        RECT 28.600 94.800 29.800 94.900 ;
        RECT 16.700 93.900 22.200 94.200 ;
        RECT 16.900 93.800 17.300 93.900 ;
        RECT 18.200 93.800 18.600 93.900 ;
        RECT 11.200 93.600 11.500 93.800 ;
        RECT 11.100 93.200 11.500 93.600 ;
        RECT 13.400 93.600 13.800 93.800 ;
        RECT 11.800 93.400 12.200 93.500 ;
        RECT 11.800 93.100 13.000 93.400 ;
        RECT 10.000 92.200 10.800 92.900 ;
        RECT 10.000 91.800 11.400 92.200 ;
        RECT 10.000 91.100 10.800 91.800 ;
        RECT 12.600 91.100 13.000 93.100 ;
        RECT 13.400 93.300 15.300 93.600 ;
        RECT 13.400 91.100 13.800 93.300 ;
        RECT 14.900 93.200 15.300 93.300 ;
        RECT 19.800 92.800 20.100 93.900 ;
        RECT 21.400 93.800 22.200 93.900 ;
        RECT 25.200 93.800 25.800 94.200 ;
        RECT 26.600 93.800 27.400 94.200 ;
        RECT 18.900 92.700 19.300 92.800 ;
        RECT 15.800 92.100 16.200 92.500 ;
        RECT 17.900 92.400 19.300 92.700 ;
        RECT 19.800 92.400 20.200 92.800 ;
        RECT 17.900 92.100 18.200 92.400 ;
        RECT 20.600 92.100 21.000 92.500 ;
        RECT 15.500 91.800 16.200 92.100 ;
        RECT 15.500 91.100 16.100 91.800 ;
        RECT 17.800 91.100 18.200 92.100 ;
        RECT 20.000 91.800 21.000 92.100 ;
        RECT 20.000 91.100 20.400 91.800 ;
        RECT 22.200 91.100 22.600 93.500 ;
        RECT 25.200 92.500 25.500 93.800 ;
        RECT 27.000 92.800 28.200 93.200 ;
        RECT 29.400 92.800 29.800 93.200 ;
        RECT 30.300 93.100 30.600 94.900 ;
        RECT 31.800 94.800 32.900 94.900 ;
        RECT 31.000 93.800 31.400 94.600 ;
        RECT 32.600 94.200 32.900 94.800 ;
        RECT 33.400 94.400 33.800 95.200 ;
        RECT 34.100 94.200 34.400 95.900 ;
        RECT 35.000 95.800 35.400 95.900 ;
        RECT 36.600 94.400 37.000 95.200 ;
        RECT 37.300 94.200 37.600 95.900 ;
        RECT 38.200 95.800 38.600 95.900 ;
        RECT 38.200 95.100 38.600 95.200 ;
        RECT 39.000 95.100 39.400 95.600 ;
        RECT 38.200 94.800 39.400 95.100 ;
        RECT 39.800 95.200 40.100 95.900 ;
        RECT 41.400 95.800 41.800 96.600 ;
        RECT 39.800 94.800 40.200 95.200 ;
        RECT 39.800 94.200 40.100 94.800 ;
        RECT 32.600 94.100 33.000 94.200 ;
        RECT 32.600 93.800 33.400 94.100 ;
        RECT 34.100 93.800 35.400 94.200 ;
        RECT 35.800 94.100 36.200 94.200 ;
        RECT 35.800 93.800 36.600 94.100 ;
        RECT 37.300 93.800 38.600 94.200 ;
        RECT 39.000 93.800 39.400 94.200 ;
        RECT 39.800 93.800 40.200 94.200 ;
        RECT 33.000 93.600 33.400 93.800 ;
        RECT 32.700 93.100 34.500 93.300 ;
        RECT 35.000 93.100 35.300 93.800 ;
        RECT 36.200 93.600 36.600 93.800 ;
        RECT 35.900 93.100 37.700 93.300 ;
        RECT 38.200 93.100 38.500 93.800 ;
        RECT 39.000 93.100 39.300 93.800 ;
        RECT 25.200 92.200 27.200 92.500 ;
        RECT 29.500 92.400 29.900 92.800 ;
        RECT 25.200 92.100 25.800 92.200 ;
        RECT 25.400 91.100 25.800 92.100 ;
        RECT 26.900 92.100 27.200 92.200 ;
        RECT 26.900 91.800 27.400 92.100 ;
        RECT 27.000 91.100 27.400 91.800 ;
        RECT 30.200 91.100 30.600 93.100 ;
        RECT 32.600 93.000 34.600 93.100 ;
        RECT 32.600 91.100 33.000 93.000 ;
        RECT 34.200 91.100 34.600 93.000 ;
        RECT 35.000 91.100 35.400 93.100 ;
        RECT 35.800 93.000 37.800 93.100 ;
        RECT 35.800 91.100 36.200 93.000 ;
        RECT 37.400 91.100 37.800 93.000 ;
        RECT 38.200 92.800 39.300 93.100 ;
        RECT 38.200 91.100 38.600 92.800 ;
        RECT 39.800 92.100 40.100 93.800 ;
        RECT 40.600 93.100 41.000 93.200 ;
        RECT 42.200 93.100 42.600 99.900 ;
        RECT 43.800 95.900 44.200 99.900 ;
        RECT 44.600 96.200 45.000 99.900 ;
        RECT 46.200 96.200 46.600 99.900 ;
        RECT 44.600 95.900 46.600 96.200 ;
        RECT 48.600 96.200 49.000 99.900 ;
        RECT 49.400 96.200 49.800 96.300 ;
        RECT 50.800 96.200 51.600 99.900 ;
        RECT 48.600 95.900 49.800 96.200 ;
        RECT 50.600 95.900 51.600 96.200 ;
        RECT 52.700 96.200 53.100 96.300 ;
        RECT 53.400 96.200 53.800 99.900 ;
        RECT 52.700 95.900 53.800 96.200 ;
        RECT 43.900 95.200 44.200 95.900 ;
        RECT 45.800 95.200 46.200 95.400 ;
        RECT 50.600 95.200 50.900 95.900 ;
        RECT 52.700 95.600 53.000 95.900 ;
        RECT 54.200 95.800 54.600 96.600 ;
        RECT 51.300 95.300 53.000 95.600 ;
        RECT 51.300 95.200 51.700 95.300 ;
        RECT 43.800 94.900 45.000 95.200 ;
        RECT 45.800 94.900 46.600 95.200 ;
        RECT 43.800 94.800 44.200 94.900 ;
        RECT 43.000 94.100 43.400 94.200 ;
        RECT 43.800 94.100 44.200 94.200 ;
        RECT 43.000 93.800 44.200 94.100 ;
        RECT 43.000 93.400 43.400 93.800 ;
        RECT 40.600 92.800 42.600 93.100 ;
        RECT 43.800 92.800 44.200 93.200 ;
        RECT 44.700 93.100 45.000 94.900 ;
        RECT 46.200 94.800 46.600 94.900 ;
        RECT 47.800 95.100 48.200 95.200 ;
        RECT 50.200 95.100 50.900 95.200 ;
        RECT 47.800 94.900 50.900 95.100 ;
        RECT 52.400 94.900 52.800 95.000 ;
        RECT 47.800 94.800 51.100 94.900 ;
        RECT 50.600 94.600 51.100 94.800 ;
        RECT 45.400 94.100 45.800 94.600 ;
        RECT 46.200 94.100 46.600 94.200 ;
        RECT 45.400 93.800 46.600 94.100 ;
        RECT 47.000 94.100 47.400 94.200 ;
        RECT 48.600 94.100 49.400 94.200 ;
        RECT 47.000 93.800 49.400 94.100 ;
        RECT 50.000 93.800 50.400 94.200 ;
        RECT 50.100 93.600 50.400 93.800 ;
        RECT 49.400 93.400 49.800 93.500 ;
        RECT 40.600 92.400 41.000 92.800 ;
        RECT 39.800 91.100 40.200 92.100 ;
        RECT 41.700 91.100 42.100 92.800 ;
        RECT 43.900 92.400 44.300 92.800 ;
        RECT 44.600 91.100 45.000 93.100 ;
        RECT 48.600 93.100 49.800 93.400 ;
        RECT 50.100 93.200 50.500 93.600 ;
        RECT 48.600 91.100 49.000 93.100 ;
        RECT 50.800 92.900 51.100 94.600 ;
        RECT 51.500 94.600 52.800 94.900 ;
        RECT 51.500 94.300 51.800 94.600 ;
        RECT 51.400 93.900 51.800 94.300 ;
        RECT 53.000 94.100 53.800 94.200 ;
        RECT 52.100 93.800 53.800 94.100 ;
        RECT 52.100 93.600 52.400 93.800 ;
        RECT 51.400 93.300 52.400 93.600 ;
        RECT 52.700 93.400 53.100 93.500 ;
        RECT 51.400 93.200 52.200 93.300 ;
        RECT 52.700 93.100 53.800 93.400 ;
        RECT 55.000 93.100 55.400 99.900 ;
        RECT 56.600 96.900 57.000 99.900 ;
        RECT 56.700 96.600 57.000 96.900 ;
        RECT 58.200 99.600 60.200 99.900 ;
        RECT 58.200 96.900 58.600 99.600 ;
        RECT 59.000 96.900 59.400 99.300 ;
        RECT 59.800 97.000 60.200 99.600 ;
        RECT 60.700 99.600 62.500 99.900 ;
        RECT 60.700 99.500 61.000 99.600 ;
        RECT 58.200 96.600 58.500 96.900 ;
        RECT 56.700 96.300 58.500 96.600 ;
        RECT 59.100 96.700 59.400 96.900 ;
        RECT 60.600 96.700 61.000 99.500 ;
        RECT 62.200 99.500 62.500 99.600 ;
        RECT 59.100 96.500 61.000 96.700 ;
        RECT 61.400 96.500 61.800 99.300 ;
        RECT 62.200 96.500 62.600 99.500 ;
        RECT 59.100 96.400 60.900 96.500 ;
        RECT 61.400 96.200 61.700 96.500 ;
        RECT 63.000 96.200 63.400 99.900 ;
        RECT 63.800 96.200 64.200 96.300 ;
        RECT 61.400 96.100 61.800 96.200 ;
        RECT 60.100 95.800 61.800 96.100 ;
        RECT 63.000 95.900 64.200 96.200 ;
        RECT 65.200 95.900 66.000 99.900 ;
        RECT 66.900 96.200 67.300 96.300 ;
        RECT 67.800 96.200 68.200 99.900 ;
        RECT 66.900 95.900 68.200 96.200 ;
        RECT 59.000 94.800 59.800 95.200 ;
        RECT 55.800 93.400 56.200 94.200 ;
        RECT 57.400 94.100 57.800 94.200 ;
        RECT 58.200 94.100 59.000 94.200 ;
        RECT 57.400 93.800 59.000 94.100 ;
        RECT 50.800 91.100 51.600 92.900 ;
        RECT 53.400 91.100 53.800 93.100 ;
        RECT 54.500 92.800 55.400 93.100 ;
        RECT 57.400 92.800 58.600 93.200 ;
        RECT 54.500 92.200 54.900 92.800 ;
        RECT 60.100 92.500 60.400 95.800 ;
        RECT 65.400 95.200 65.700 95.900 ;
        RECT 66.300 95.200 66.700 95.300 ;
        RECT 61.400 95.100 61.800 95.200 ;
        RECT 65.400 95.100 65.800 95.200 ;
        RECT 61.400 94.800 65.800 95.100 ;
        RECT 66.300 94.900 67.100 95.200 ;
        RECT 66.700 94.800 67.100 94.900 ;
        RECT 65.400 94.200 65.700 94.800 ;
        RECT 63.000 93.800 63.800 94.200 ;
        RECT 64.400 93.800 64.800 94.200 ;
        RECT 64.500 93.600 64.800 93.800 ;
        RECT 65.200 93.900 65.700 94.200 ;
        RECT 66.000 94.300 66.400 94.400 ;
        RECT 66.000 94.200 67.400 94.300 ;
        RECT 66.000 94.000 68.200 94.200 ;
        RECT 67.100 93.900 68.200 94.000 ;
        RECT 63.800 93.400 64.200 93.500 ;
        RECT 58.400 92.200 60.400 92.500 ;
        RECT 54.200 91.800 54.900 92.200 ;
        RECT 54.500 91.100 54.900 91.800 ;
        RECT 58.200 91.800 58.700 92.200 ;
        RECT 59.800 92.100 60.400 92.200 ;
        RECT 63.000 93.100 64.200 93.400 ;
        RECT 64.500 93.200 64.900 93.600 ;
        RECT 58.200 91.100 58.600 91.800 ;
        RECT 59.800 91.100 60.200 92.100 ;
        RECT 63.000 91.100 63.400 93.100 ;
        RECT 65.200 92.900 65.500 93.900 ;
        RECT 67.400 93.800 68.200 93.900 ;
        RECT 69.400 94.100 69.800 99.900 ;
        RECT 71.500 96.200 71.900 99.900 ;
        RECT 73.400 97.500 73.800 99.500 ;
        RECT 72.200 96.800 72.600 97.200 ;
        RECT 72.300 96.200 72.600 96.800 ;
        RECT 71.500 95.900 72.000 96.200 ;
        RECT 72.300 95.900 73.000 96.200 ;
        RECT 71.000 94.400 71.400 95.200 ;
        RECT 71.700 94.200 72.000 95.900 ;
        RECT 72.600 95.800 73.000 95.900 ;
        RECT 73.400 95.800 73.700 97.500 ;
        RECT 75.500 96.400 75.900 99.900 ;
        RECT 75.500 96.100 76.300 96.400 ;
        RECT 73.400 95.500 75.300 95.800 ;
        RECT 73.400 94.400 73.800 95.200 ;
        RECT 74.200 94.400 74.600 95.200 ;
        RECT 75.000 94.500 75.300 95.500 ;
        RECT 70.200 94.100 70.600 94.200 ;
        RECT 69.400 93.800 71.000 94.100 ;
        RECT 71.700 93.800 73.000 94.200 ;
        RECT 75.000 94.100 75.700 94.500 ;
        RECT 76.000 94.200 76.300 96.100 ;
        RECT 78.500 96.300 78.900 99.900 ;
        RECT 80.600 97.500 81.000 99.500 ;
        RECT 78.500 95.900 79.400 96.300 ;
        RECT 76.600 95.100 77.000 95.600 ;
        RECT 77.400 95.100 77.800 95.200 ;
        RECT 76.600 94.800 77.800 95.100 ;
        RECT 78.200 94.800 78.600 95.600 ;
        RECT 76.000 94.100 77.000 94.200 ;
        RECT 78.200 94.100 78.500 94.800 ;
        RECT 75.000 93.900 75.500 94.100 ;
        RECT 65.800 93.200 66.600 93.600 ;
        RECT 66.900 93.400 67.300 93.500 ;
        RECT 66.900 93.100 68.200 93.400 ;
        RECT 65.200 91.100 66.000 92.900 ;
        RECT 67.800 91.100 68.200 93.100 ;
        RECT 68.600 92.400 69.000 93.200 ;
        RECT 69.400 91.100 69.800 93.800 ;
        RECT 70.600 93.600 71.000 93.800 ;
        RECT 70.300 93.100 72.100 93.300 ;
        RECT 72.600 93.100 72.900 93.800 ;
        RECT 73.400 93.600 75.500 93.900 ;
        RECT 76.000 93.800 78.500 94.100 ;
        RECT 79.000 94.200 79.300 95.900 ;
        RECT 80.600 95.800 80.900 97.500 ;
        RECT 82.700 96.400 83.100 99.900 ;
        RECT 82.700 96.100 83.500 96.400 ;
        RECT 80.600 95.500 82.500 95.800 ;
        RECT 80.600 94.400 81.000 95.200 ;
        RECT 81.400 94.400 81.800 95.200 ;
        RECT 82.200 94.500 82.500 95.500 ;
        RECT 79.000 93.800 79.400 94.200 ;
        RECT 82.200 94.100 82.900 94.500 ;
        RECT 83.200 94.200 83.500 96.100 ;
        RECT 85.700 96.300 86.100 99.900 ;
        RECT 85.700 95.900 86.600 96.300 ;
        RECT 83.800 94.800 84.200 95.600 ;
        RECT 85.400 94.800 85.800 95.600 ;
        RECT 83.200 94.100 84.200 94.200 ;
        RECT 85.400 94.100 85.700 94.800 ;
        RECT 82.200 93.900 82.700 94.100 ;
        RECT 70.200 93.000 72.200 93.100 ;
        RECT 70.200 91.100 70.600 93.000 ;
        RECT 71.800 91.100 72.200 93.000 ;
        RECT 72.600 91.100 73.000 93.100 ;
        RECT 73.400 92.500 73.700 93.600 ;
        RECT 76.000 93.500 76.300 93.800 ;
        RECT 75.900 93.300 76.300 93.500 ;
        RECT 75.500 93.000 76.300 93.300 ;
        RECT 73.400 91.500 73.800 92.500 ;
        RECT 75.500 91.500 75.900 93.000 ;
        RECT 79.000 92.200 79.300 93.800 ;
        RECT 80.600 93.600 82.700 93.900 ;
        RECT 83.200 93.800 85.700 94.100 ;
        RECT 86.200 94.200 86.500 95.900 ;
        RECT 87.800 95.600 88.200 99.900 ;
        RECT 89.900 97.900 90.500 99.900 ;
        RECT 92.200 97.900 92.600 99.900 ;
        RECT 94.400 98.200 94.800 99.900 ;
        RECT 94.400 97.900 95.400 98.200 ;
        RECT 90.200 97.500 90.600 97.900 ;
        RECT 92.300 97.600 92.600 97.900 ;
        RECT 91.900 97.300 93.700 97.600 ;
        RECT 95.000 97.500 95.400 97.900 ;
        RECT 91.900 97.200 92.300 97.300 ;
        RECT 93.300 97.200 93.700 97.300 ;
        RECT 89.800 96.600 90.500 97.000 ;
        RECT 90.200 96.100 90.500 96.600 ;
        RECT 91.300 96.500 92.400 96.800 ;
        RECT 91.300 96.400 91.700 96.500 ;
        RECT 90.200 95.800 91.400 96.100 ;
        RECT 87.800 95.300 89.900 95.600 ;
        RECT 87.000 94.800 87.400 95.200 ;
        RECT 86.200 94.100 86.600 94.200 ;
        RECT 87.000 94.100 87.300 94.800 ;
        RECT 86.200 93.800 87.300 94.100 ;
        RECT 79.800 92.400 80.200 93.200 ;
        RECT 80.600 92.500 80.900 93.600 ;
        RECT 83.200 93.500 83.500 93.800 ;
        RECT 83.100 93.300 83.500 93.500 ;
        RECT 82.700 93.000 83.500 93.300 ;
        RECT 79.000 91.100 79.400 92.200 ;
        RECT 80.600 91.500 81.000 92.500 ;
        RECT 82.700 91.500 83.100 93.000 ;
        RECT 86.200 92.100 86.500 93.800 ;
        RECT 87.800 93.600 88.200 95.300 ;
        RECT 89.500 95.200 89.900 95.300 ;
        RECT 91.100 95.200 91.400 95.800 ;
        RECT 92.100 95.900 92.400 96.500 ;
        RECT 92.700 96.500 93.100 96.600 ;
        RECT 95.000 96.500 95.400 96.600 ;
        RECT 92.700 96.200 95.400 96.500 ;
        RECT 92.100 95.700 94.500 95.900 ;
        RECT 96.600 95.700 97.000 99.900 ;
        RECT 92.100 95.600 97.000 95.700 ;
        RECT 94.100 95.500 97.000 95.600 ;
        RECT 94.200 95.400 97.000 95.500 ;
        RECT 99.800 95.600 100.200 99.900 ;
        RECT 101.400 95.600 101.800 99.900 ;
        RECT 103.000 95.600 103.400 99.900 ;
        RECT 104.600 95.600 105.000 99.900 ;
        RECT 107.500 96.300 107.900 99.900 ;
        RECT 107.000 95.900 107.900 96.300 ;
        RECT 108.600 97.500 109.000 99.500 ;
        RECT 99.800 95.200 100.700 95.600 ;
        RECT 101.400 95.200 102.500 95.600 ;
        RECT 103.000 95.200 104.100 95.600 ;
        RECT 104.600 95.200 105.800 95.600 ;
        RECT 88.700 94.900 89.100 95.000 ;
        RECT 88.700 94.600 90.600 94.900 ;
        RECT 91.000 94.800 91.400 95.200 ;
        RECT 93.400 95.100 93.800 95.200 ;
        RECT 93.400 94.800 95.900 95.100 ;
        RECT 90.200 94.500 90.600 94.600 ;
        RECT 91.100 94.200 91.400 94.800 ;
        RECT 95.500 94.700 95.900 94.800 ;
        RECT 100.300 94.500 100.700 95.200 ;
        RECT 102.100 94.500 102.500 95.200 ;
        RECT 103.700 94.500 104.100 95.200 ;
        RECT 94.700 94.200 95.100 94.300 ;
        RECT 91.100 93.900 96.600 94.200 ;
        RECT 91.300 93.800 91.700 93.900 ;
        RECT 87.800 93.300 89.700 93.600 ;
        RECT 87.000 92.400 87.400 93.200 ;
        RECT 86.200 91.100 86.600 92.100 ;
        RECT 87.800 91.100 88.200 93.300 ;
        RECT 89.300 93.200 89.700 93.300 ;
        RECT 94.200 92.800 94.500 93.900 ;
        RECT 95.800 93.800 96.600 93.900 ;
        RECT 100.300 94.100 101.600 94.500 ;
        RECT 102.100 94.100 103.300 94.500 ;
        RECT 103.700 94.100 105.000 94.500 ;
        RECT 100.300 93.800 100.700 94.100 ;
        RECT 102.100 93.800 102.500 94.100 ;
        RECT 103.700 93.800 104.100 94.100 ;
        RECT 105.400 93.800 105.800 95.200 ;
        RECT 107.100 94.200 107.400 95.900 ;
        RECT 108.600 95.800 108.900 97.500 ;
        RECT 110.700 96.400 111.100 99.900 ;
        RECT 113.800 96.800 114.200 97.200 ;
        RECT 110.700 96.100 111.500 96.400 ;
        RECT 113.800 96.200 114.100 96.800 ;
        RECT 114.500 96.200 114.900 99.900 ;
        RECT 107.800 94.800 108.200 95.600 ;
        RECT 108.600 95.500 110.500 95.800 ;
        RECT 108.600 94.400 109.000 95.200 ;
        RECT 109.400 94.400 109.800 95.200 ;
        RECT 110.200 94.500 110.500 95.500 ;
        RECT 107.000 93.800 107.400 94.200 ;
        RECT 110.200 94.100 110.900 94.500 ;
        RECT 111.200 94.200 111.500 96.100 ;
        RECT 113.400 95.900 114.100 96.200 ;
        RECT 114.400 95.900 114.900 96.200 ;
        RECT 113.400 95.800 113.800 95.900 ;
        RECT 111.800 94.800 112.200 95.600 ;
        RECT 114.400 94.200 114.700 95.900 ;
        RECT 116.600 95.800 117.000 96.600 ;
        RECT 115.000 95.100 115.400 95.200 ;
        RECT 116.600 95.100 116.900 95.800 ;
        RECT 115.000 94.800 116.900 95.100 ;
        RECT 115.000 94.400 115.400 94.800 ;
        RECT 110.200 93.900 110.700 94.100 ;
        RECT 93.300 92.700 93.700 92.800 ;
        RECT 90.200 92.100 90.600 92.500 ;
        RECT 92.300 92.400 93.700 92.700 ;
        RECT 94.200 92.400 94.600 92.800 ;
        RECT 92.300 92.100 92.600 92.400 ;
        RECT 95.000 92.100 95.400 92.500 ;
        RECT 89.900 91.800 90.600 92.100 ;
        RECT 89.900 91.100 90.500 91.800 ;
        RECT 92.200 91.100 92.600 92.100 ;
        RECT 94.400 91.800 95.400 92.100 ;
        RECT 94.400 91.100 94.800 91.800 ;
        RECT 96.600 91.100 97.000 93.500 ;
        RECT 99.800 93.400 100.700 93.800 ;
        RECT 101.400 93.400 102.500 93.800 ;
        RECT 103.000 93.400 104.100 93.800 ;
        RECT 104.600 93.400 105.800 93.800 ;
        RECT 99.800 91.100 100.200 93.400 ;
        RECT 101.400 91.100 101.800 93.400 ;
        RECT 103.000 91.100 103.400 93.400 ;
        RECT 104.600 91.100 105.000 93.400 ;
        RECT 106.200 92.400 106.600 93.200 ;
        RECT 107.100 92.200 107.400 93.800 ;
        RECT 107.000 91.100 107.400 92.200 ;
        RECT 108.600 93.600 110.700 93.900 ;
        RECT 111.200 93.800 112.200 94.200 ;
        RECT 113.400 93.800 114.700 94.200 ;
        RECT 115.800 94.100 116.200 94.200 ;
        RECT 115.400 93.800 116.200 94.100 ;
        RECT 116.600 94.100 117.000 94.200 ;
        RECT 117.400 94.100 117.800 99.900 ;
        RECT 116.600 93.800 117.800 94.100 ;
        RECT 108.600 92.500 108.900 93.600 ;
        RECT 111.200 93.500 111.500 93.800 ;
        RECT 111.100 93.300 111.500 93.500 ;
        RECT 110.700 93.200 111.500 93.300 ;
        RECT 110.200 93.000 111.500 93.200 ;
        RECT 113.500 93.100 113.800 93.800 ;
        RECT 115.400 93.600 115.800 93.800 ;
        RECT 114.300 93.100 116.100 93.300 ;
        RECT 117.400 93.100 117.800 93.800 ;
        RECT 118.200 93.400 118.600 94.200 ;
        RECT 110.200 92.800 111.100 93.000 ;
        RECT 108.600 91.500 109.000 92.500 ;
        RECT 110.700 91.500 111.100 92.800 ;
        RECT 113.400 91.100 113.800 93.100 ;
        RECT 114.200 93.000 116.200 93.100 ;
        RECT 114.200 91.100 114.600 93.000 ;
        RECT 115.800 91.100 116.200 93.000 ;
        RECT 116.900 92.800 117.800 93.100 ;
        RECT 116.900 91.100 117.300 92.800 ;
        RECT 119.000 91.100 119.400 99.900 ;
        RECT 121.000 96.800 121.400 97.200 ;
        RECT 121.000 96.200 121.300 96.800 ;
        RECT 121.700 96.200 122.100 99.900 ;
        RECT 120.600 95.900 121.300 96.200 ;
        RECT 121.600 95.900 122.100 96.200 ;
        RECT 120.600 95.800 121.000 95.900 ;
        RECT 121.600 94.200 121.900 95.900 ;
        RECT 122.200 94.400 122.600 95.200 ;
        RECT 120.600 93.800 121.900 94.200 ;
        RECT 123.000 94.100 123.400 94.200 ;
        RECT 123.800 94.100 124.200 99.900 ;
        RECT 125.400 96.200 125.800 99.900 ;
        RECT 126.200 96.200 126.600 96.300 ;
        RECT 125.400 95.900 126.600 96.200 ;
        RECT 127.600 95.900 128.400 99.900 ;
        RECT 129.300 96.200 129.700 96.300 ;
        RECT 130.200 96.200 130.600 99.900 ;
        RECT 131.000 96.900 131.400 99.900 ;
        RECT 131.100 96.600 131.400 96.900 ;
        RECT 132.600 99.600 134.600 99.900 ;
        RECT 132.600 96.900 133.000 99.600 ;
        RECT 133.400 96.900 133.800 99.300 ;
        RECT 134.200 97.000 134.600 99.600 ;
        RECT 135.100 99.600 136.900 99.900 ;
        RECT 135.100 99.500 135.400 99.600 ;
        RECT 132.600 96.600 132.900 96.900 ;
        RECT 131.100 96.300 132.900 96.600 ;
        RECT 133.500 96.700 133.800 96.900 ;
        RECT 135.000 96.700 135.400 99.500 ;
        RECT 136.600 99.500 136.900 99.600 ;
        RECT 133.500 96.500 135.400 96.700 ;
        RECT 135.800 96.500 136.200 99.300 ;
        RECT 136.600 96.500 137.000 99.500 ;
        RECT 133.500 96.400 135.300 96.500 ;
        RECT 129.300 95.900 130.600 96.200 ;
        RECT 135.800 96.200 136.100 96.500 ;
        RECT 137.400 96.200 137.800 99.900 ;
        RECT 138.300 96.200 138.700 96.300 ;
        RECT 135.800 96.100 136.200 96.200 ;
        RECT 127.800 95.200 128.100 95.900 ;
        RECT 134.500 95.800 136.200 96.100 ;
        RECT 137.400 95.900 138.700 96.200 ;
        RECT 139.600 95.900 140.400 99.900 ;
        RECT 141.400 96.200 141.800 96.300 ;
        RECT 142.200 96.200 142.600 99.900 ;
        RECT 141.400 95.900 142.600 96.200 ;
        RECT 128.700 95.200 129.100 95.300 ;
        RECT 127.800 94.800 128.200 95.200 ;
        RECT 128.700 94.900 129.500 95.200 ;
        RECT 129.100 94.800 129.500 94.900 ;
        RECT 133.400 94.800 134.200 95.200 ;
        RECT 127.800 94.200 128.100 94.800 ;
        RECT 122.600 93.800 124.200 94.100 ;
        RECT 125.400 93.800 126.200 94.200 ;
        RECT 126.800 93.800 127.200 94.200 ;
        RECT 119.800 92.400 120.200 93.200 ;
        RECT 120.700 93.100 121.000 93.800 ;
        RECT 122.600 93.600 123.000 93.800 ;
        RECT 121.500 93.100 123.300 93.300 ;
        RECT 120.600 91.100 121.000 93.100 ;
        RECT 121.400 93.000 123.400 93.100 ;
        RECT 121.400 91.100 121.800 93.000 ;
        RECT 123.000 91.100 123.400 93.000 ;
        RECT 123.800 91.100 124.200 93.800 ;
        RECT 126.900 93.600 127.200 93.800 ;
        RECT 127.600 93.900 128.100 94.200 ;
        RECT 128.400 94.300 128.800 94.400 ;
        RECT 128.400 94.200 129.800 94.300 ;
        RECT 128.400 94.000 130.600 94.200 ;
        RECT 129.500 93.900 130.600 94.000 ;
        RECT 126.200 93.400 126.600 93.500 ;
        RECT 124.600 92.400 125.000 93.200 ;
        RECT 125.400 93.100 126.600 93.400 ;
        RECT 126.900 93.200 127.300 93.600 ;
        RECT 125.400 91.100 125.800 93.100 ;
        RECT 127.600 92.900 127.900 93.900 ;
        RECT 129.800 93.800 130.600 93.900 ;
        RECT 132.600 93.800 133.800 94.200 ;
        RECT 128.200 93.200 129.000 93.600 ;
        RECT 129.300 93.400 129.700 93.500 ;
        RECT 129.300 93.100 130.600 93.400 ;
        RECT 127.600 92.200 128.400 92.900 ;
        RECT 127.600 91.800 129.000 92.200 ;
        RECT 127.600 91.100 128.400 91.800 ;
        RECT 130.200 91.100 130.600 93.100 ;
        RECT 131.000 93.100 131.400 93.200 ;
        RECT 131.800 93.100 132.700 93.200 ;
        RECT 131.000 92.800 132.700 93.100 ;
        RECT 134.500 92.500 134.800 95.800 ;
        RECT 138.900 95.200 139.300 95.300 ;
        RECT 139.900 95.200 140.200 95.900 ;
        RECT 138.500 94.900 139.300 95.200 ;
        RECT 138.500 94.800 138.900 94.900 ;
        RECT 139.800 94.800 140.200 95.200 ;
        RECT 139.200 94.300 139.600 94.400 ;
        RECT 138.200 94.200 139.600 94.300 ;
        RECT 137.400 94.000 139.600 94.200 ;
        RECT 139.900 94.200 140.200 94.800 ;
        RECT 143.000 95.600 143.400 99.900 ;
        RECT 145.100 97.900 145.700 99.900 ;
        RECT 147.400 97.900 147.800 99.900 ;
        RECT 149.600 98.200 150.000 99.900 ;
        RECT 149.600 97.900 150.600 98.200 ;
        RECT 145.400 97.500 145.800 97.900 ;
        RECT 147.500 97.600 147.800 97.900 ;
        RECT 147.100 97.300 148.900 97.600 ;
        RECT 150.200 97.500 150.600 97.900 ;
        RECT 147.100 97.200 147.500 97.300 ;
        RECT 148.500 97.200 148.900 97.300 ;
        RECT 145.000 96.600 145.700 97.000 ;
        RECT 145.400 96.100 145.700 96.600 ;
        RECT 146.500 96.500 147.600 96.800 ;
        RECT 146.500 96.400 146.900 96.500 ;
        RECT 145.400 95.800 146.600 96.100 ;
        RECT 143.000 95.300 145.100 95.600 ;
        RECT 137.400 93.900 138.500 94.000 ;
        RECT 139.900 93.900 140.400 94.200 ;
        RECT 137.400 93.800 138.200 93.900 ;
        RECT 138.300 93.400 138.700 93.500 ;
        RECT 132.800 92.200 134.800 92.500 ;
        RECT 132.600 91.800 133.100 92.200 ;
        RECT 134.200 92.100 134.800 92.200 ;
        RECT 137.400 93.100 138.700 93.400 ;
        RECT 139.000 93.200 139.800 93.600 ;
        RECT 132.600 91.100 133.000 91.800 ;
        RECT 134.200 91.100 134.600 92.100 ;
        RECT 137.400 91.100 137.800 93.100 ;
        RECT 140.100 92.900 140.400 93.900 ;
        RECT 140.800 93.800 141.200 94.200 ;
        RECT 141.800 93.800 142.600 94.200 ;
        RECT 140.800 93.600 141.100 93.800 ;
        RECT 140.700 93.200 141.100 93.600 ;
        RECT 143.000 93.600 143.400 95.300 ;
        RECT 144.700 95.200 145.100 95.300 ;
        RECT 143.900 94.900 144.300 95.000 ;
        RECT 143.900 94.600 145.800 94.900 ;
        RECT 145.400 94.500 145.800 94.600 ;
        RECT 146.300 94.200 146.600 95.800 ;
        RECT 147.300 95.900 147.600 96.500 ;
        RECT 147.900 96.500 148.300 96.600 ;
        RECT 150.200 96.500 150.600 96.600 ;
        RECT 147.900 96.200 150.600 96.500 ;
        RECT 147.300 95.700 149.700 95.900 ;
        RECT 151.800 95.700 152.200 99.900 ;
        RECT 147.300 95.600 152.200 95.700 ;
        RECT 149.300 95.500 152.200 95.600 ;
        RECT 149.400 95.400 152.200 95.500 ;
        RECT 154.200 95.600 154.600 99.900 ;
        RECT 156.300 97.900 156.900 99.900 ;
        RECT 158.600 97.900 159.000 99.900 ;
        RECT 160.800 98.200 161.200 99.900 ;
        RECT 160.800 97.900 161.800 98.200 ;
        RECT 156.600 97.500 157.000 97.900 ;
        RECT 158.700 97.600 159.000 97.900 ;
        RECT 158.300 97.300 160.100 97.600 ;
        RECT 161.400 97.500 161.800 97.900 ;
        RECT 158.300 97.200 158.700 97.300 ;
        RECT 159.700 97.200 160.100 97.300 ;
        RECT 156.200 96.600 156.900 97.000 ;
        RECT 156.600 96.100 156.900 96.600 ;
        RECT 157.700 96.500 158.800 96.800 ;
        RECT 157.700 96.400 158.100 96.500 ;
        RECT 156.600 95.800 157.800 96.100 ;
        RECT 154.200 95.300 156.300 95.600 ;
        RECT 148.600 95.100 149.000 95.200 ;
        RECT 148.600 94.800 151.100 95.100 ;
        RECT 149.400 94.700 149.800 94.800 ;
        RECT 150.700 94.700 151.100 94.800 ;
        RECT 149.900 94.200 150.300 94.300 ;
        RECT 146.300 93.900 151.800 94.200 ;
        RECT 146.500 93.800 146.900 93.900 ;
        RECT 141.400 93.400 141.800 93.500 ;
        RECT 141.400 93.100 142.600 93.400 ;
        RECT 139.600 92.200 140.400 92.900 ;
        RECT 139.000 91.800 140.400 92.200 ;
        RECT 139.600 91.100 140.400 91.800 ;
        RECT 142.200 91.100 142.600 93.100 ;
        RECT 143.000 93.300 144.900 93.600 ;
        RECT 143.000 91.100 143.400 93.300 ;
        RECT 144.500 93.200 144.900 93.300 ;
        RECT 149.400 92.800 149.700 93.900 ;
        RECT 151.000 93.800 151.800 93.900 ;
        RECT 154.200 93.600 154.600 95.300 ;
        RECT 155.900 95.200 156.300 95.300 ;
        RECT 155.100 94.900 155.500 95.000 ;
        RECT 155.100 94.600 157.000 94.900 ;
        RECT 156.600 94.500 157.000 94.600 ;
        RECT 157.500 94.200 157.800 95.800 ;
        RECT 158.500 95.900 158.800 96.500 ;
        RECT 159.100 96.500 159.500 96.600 ;
        RECT 161.400 96.500 161.800 96.600 ;
        RECT 159.100 96.200 161.800 96.500 ;
        RECT 158.500 95.700 160.900 95.900 ;
        RECT 163.000 95.700 163.400 99.900 ;
        RECT 158.500 95.600 163.400 95.700 ;
        RECT 160.500 95.500 163.400 95.600 ;
        RECT 160.600 95.400 163.400 95.500 ;
        RECT 163.800 95.700 164.200 99.900 ;
        RECT 166.000 98.200 166.400 99.900 ;
        RECT 165.400 97.900 166.400 98.200 ;
        RECT 168.200 97.900 168.600 99.900 ;
        RECT 170.300 97.900 170.900 99.900 ;
        RECT 165.400 97.500 165.800 97.900 ;
        RECT 168.200 97.600 168.500 97.900 ;
        RECT 167.100 97.300 168.900 97.600 ;
        RECT 170.200 97.500 170.600 97.900 ;
        RECT 167.100 97.200 167.500 97.300 ;
        RECT 168.500 97.200 168.900 97.300 ;
        RECT 165.400 96.500 165.800 96.600 ;
        RECT 167.700 96.500 168.100 96.600 ;
        RECT 165.400 96.200 168.100 96.500 ;
        RECT 168.400 96.500 169.500 96.800 ;
        RECT 168.400 95.900 168.700 96.500 ;
        RECT 169.100 96.400 169.500 96.500 ;
        RECT 170.300 96.600 171.000 97.000 ;
        RECT 170.300 96.100 170.600 96.600 ;
        RECT 166.300 95.700 168.700 95.900 ;
        RECT 163.800 95.600 168.700 95.700 ;
        RECT 169.400 95.800 170.600 96.100 ;
        RECT 163.800 95.500 166.700 95.600 ;
        RECT 163.800 95.400 166.600 95.500 ;
        RECT 169.400 95.200 169.700 95.800 ;
        RECT 172.600 95.600 173.000 99.900 ;
        RECT 170.900 95.300 173.000 95.600 ;
        RECT 170.900 95.200 171.300 95.300 ;
        RECT 159.800 95.100 160.200 95.200 ;
        RECT 167.000 95.100 167.400 95.200 ;
        RECT 159.800 94.800 162.300 95.100 ;
        RECT 161.900 94.700 162.300 94.800 ;
        RECT 164.900 94.800 167.400 95.100 ;
        RECT 169.400 94.800 169.800 95.200 ;
        RECT 171.700 94.900 172.100 95.000 ;
        RECT 164.900 94.700 165.300 94.800 ;
        RECT 166.200 94.700 166.600 94.800 ;
        RECT 161.100 94.200 161.500 94.300 ;
        RECT 165.700 94.200 166.100 94.300 ;
        RECT 169.400 94.200 169.700 94.800 ;
        RECT 170.200 94.600 172.100 94.900 ;
        RECT 170.200 94.500 170.600 94.600 ;
        RECT 157.500 94.100 163.000 94.200 ;
        RECT 164.200 94.100 169.700 94.200 ;
        RECT 157.500 93.900 169.700 94.100 ;
        RECT 157.700 93.800 158.100 93.900 ;
        RECT 148.500 92.700 148.900 92.800 ;
        RECT 145.400 92.100 145.800 92.500 ;
        RECT 147.500 92.400 148.900 92.700 ;
        RECT 149.400 92.400 149.800 92.800 ;
        RECT 147.500 92.100 147.800 92.400 ;
        RECT 150.200 92.100 150.600 92.500 ;
        RECT 145.100 91.800 145.800 92.100 ;
        RECT 145.100 91.100 145.700 91.800 ;
        RECT 147.400 91.100 147.800 92.100 ;
        RECT 149.600 91.800 150.600 92.100 ;
        RECT 149.600 91.100 150.000 91.800 ;
        RECT 151.800 91.100 152.200 93.500 ;
        RECT 154.200 93.300 156.100 93.600 ;
        RECT 154.200 91.100 154.600 93.300 ;
        RECT 155.700 93.200 156.100 93.300 ;
        RECT 160.600 92.800 160.900 93.900 ;
        RECT 162.200 93.800 165.000 93.900 ;
        RECT 159.700 92.700 160.100 92.800 ;
        RECT 156.600 92.100 157.000 92.500 ;
        RECT 158.700 92.400 160.100 92.700 ;
        RECT 160.600 92.400 161.000 92.800 ;
        RECT 158.700 92.100 159.000 92.400 ;
        RECT 161.400 92.100 161.800 92.500 ;
        RECT 156.300 91.800 157.000 92.100 ;
        RECT 156.300 91.100 156.900 91.800 ;
        RECT 158.600 91.100 159.000 92.100 ;
        RECT 160.800 91.800 161.800 92.100 ;
        RECT 160.800 91.100 161.200 91.800 ;
        RECT 163.000 91.100 163.400 93.500 ;
        RECT 163.800 91.100 164.200 93.500 ;
        RECT 166.300 92.800 166.600 93.900 ;
        RECT 169.100 93.800 169.500 93.900 ;
        RECT 172.600 93.600 173.000 95.300 ;
        RECT 171.100 93.300 173.000 93.600 ;
        RECT 171.100 93.200 171.500 93.300 ;
        RECT 165.400 92.100 165.800 92.500 ;
        RECT 166.200 92.400 166.600 92.800 ;
        RECT 167.100 92.700 167.500 92.800 ;
        RECT 167.100 92.400 168.500 92.700 ;
        RECT 168.200 92.100 168.500 92.400 ;
        RECT 170.200 92.100 170.600 92.500 ;
        RECT 165.400 91.800 166.400 92.100 ;
        RECT 166.000 91.100 166.400 91.800 ;
        RECT 168.200 91.100 168.600 92.100 ;
        RECT 170.200 91.800 170.900 92.100 ;
        RECT 170.300 91.100 170.900 91.800 ;
        RECT 172.600 91.100 173.000 93.300 ;
        RECT 173.400 95.600 173.800 99.900 ;
        RECT 175.500 97.900 176.100 99.900 ;
        RECT 177.800 97.900 178.200 99.900 ;
        RECT 180.000 98.200 180.400 99.900 ;
        RECT 180.000 97.900 181.000 98.200 ;
        RECT 175.800 97.500 176.200 97.900 ;
        RECT 177.900 97.600 178.200 97.900 ;
        RECT 177.500 97.300 179.300 97.600 ;
        RECT 180.600 97.500 181.000 97.900 ;
        RECT 177.500 97.200 177.900 97.300 ;
        RECT 178.900 97.200 179.300 97.300 ;
        RECT 175.400 96.600 176.100 97.000 ;
        RECT 175.800 96.100 176.100 96.600 ;
        RECT 176.900 96.500 178.000 96.800 ;
        RECT 176.900 96.400 177.300 96.500 ;
        RECT 175.800 95.800 177.000 96.100 ;
        RECT 173.400 95.300 175.500 95.600 ;
        RECT 173.400 93.600 173.800 95.300 ;
        RECT 175.100 95.200 175.500 95.300 ;
        RECT 176.700 95.200 177.000 95.800 ;
        RECT 177.700 95.900 178.000 96.500 ;
        RECT 178.300 96.500 178.700 96.600 ;
        RECT 180.600 96.500 181.000 96.600 ;
        RECT 178.300 96.200 181.000 96.500 ;
        RECT 177.700 95.700 180.100 95.900 ;
        RECT 182.200 95.700 182.600 99.900 ;
        RECT 177.700 95.600 182.600 95.700 ;
        RECT 179.700 95.500 182.600 95.600 ;
        RECT 179.800 95.400 182.600 95.500 ;
        RECT 183.000 95.700 183.400 99.900 ;
        RECT 185.200 98.200 185.600 99.900 ;
        RECT 184.600 97.900 185.600 98.200 ;
        RECT 187.400 97.900 187.800 99.900 ;
        RECT 189.500 97.900 190.100 99.900 ;
        RECT 184.600 97.500 185.000 97.900 ;
        RECT 187.400 97.600 187.700 97.900 ;
        RECT 186.300 97.300 188.100 97.600 ;
        RECT 189.400 97.500 189.800 97.900 ;
        RECT 186.300 97.200 186.700 97.300 ;
        RECT 187.700 97.200 188.100 97.300 ;
        RECT 184.600 96.500 185.000 96.600 ;
        RECT 186.900 96.500 187.300 96.600 ;
        RECT 184.600 96.200 187.300 96.500 ;
        RECT 187.600 96.500 188.700 96.800 ;
        RECT 187.600 95.900 187.900 96.500 ;
        RECT 188.300 96.400 188.700 96.500 ;
        RECT 189.500 96.600 190.200 97.000 ;
        RECT 189.500 96.100 189.800 96.600 ;
        RECT 185.500 95.700 187.900 95.900 ;
        RECT 183.000 95.600 187.900 95.700 ;
        RECT 188.600 95.800 189.800 96.100 ;
        RECT 183.000 95.500 185.900 95.600 ;
        RECT 183.000 95.400 185.800 95.500 ;
        RECT 174.300 94.900 174.700 95.000 ;
        RECT 174.300 94.600 176.200 94.900 ;
        RECT 176.600 94.800 177.000 95.200 ;
        RECT 179.000 95.100 179.400 95.200 ;
        RECT 186.200 95.100 186.600 95.200 ;
        RECT 179.000 94.800 181.500 95.100 ;
        RECT 175.800 94.500 176.200 94.600 ;
        RECT 176.700 94.200 177.000 94.800 ;
        RECT 181.100 94.700 181.500 94.800 ;
        RECT 184.100 94.800 186.600 95.100 ;
        RECT 184.100 94.700 184.500 94.800 ;
        RECT 185.400 94.700 185.800 94.800 ;
        RECT 180.300 94.200 180.700 94.300 ;
        RECT 184.900 94.200 185.300 94.300 ;
        RECT 188.600 94.200 188.900 95.800 ;
        RECT 191.800 95.600 192.200 99.900 ;
        RECT 192.600 96.200 193.000 99.900 ;
        RECT 192.600 95.900 193.700 96.200 ;
        RECT 190.100 95.300 192.200 95.600 ;
        RECT 190.100 95.200 190.500 95.300 ;
        RECT 190.900 94.900 191.300 95.000 ;
        RECT 189.400 94.600 191.300 94.900 ;
        RECT 189.400 94.500 189.800 94.600 ;
        RECT 176.700 93.900 182.200 94.200 ;
        RECT 176.900 93.800 177.300 93.900 ;
        RECT 173.400 93.300 175.300 93.600 ;
        RECT 173.400 91.100 173.800 93.300 ;
        RECT 174.900 93.200 175.300 93.300 ;
        RECT 179.800 92.800 180.100 93.900 ;
        RECT 181.400 93.800 182.200 93.900 ;
        RECT 183.400 93.900 188.900 94.200 ;
        RECT 183.400 93.800 184.200 93.900 ;
        RECT 178.900 92.700 179.300 92.800 ;
        RECT 175.800 92.100 176.200 92.500 ;
        RECT 177.900 92.400 179.300 92.700 ;
        RECT 179.800 92.400 180.200 92.800 ;
        RECT 177.900 92.100 178.200 92.400 ;
        RECT 180.600 92.100 181.000 92.500 ;
        RECT 175.500 91.800 176.200 92.100 ;
        RECT 175.500 91.100 176.100 91.800 ;
        RECT 177.800 91.100 178.200 92.100 ;
        RECT 180.000 91.800 181.000 92.100 ;
        RECT 180.000 91.100 180.400 91.800 ;
        RECT 182.200 91.100 182.600 93.500 ;
        RECT 183.000 91.100 183.400 93.500 ;
        RECT 185.500 92.800 185.800 93.900 ;
        RECT 188.300 93.800 188.700 93.900 ;
        RECT 191.800 93.600 192.200 95.300 ;
        RECT 193.400 95.600 193.700 95.900 ;
        RECT 193.400 95.200 194.000 95.600 ;
        RECT 193.400 93.700 193.700 95.200 ;
        RECT 190.300 93.300 192.200 93.600 ;
        RECT 190.300 93.200 190.700 93.300 ;
        RECT 184.600 92.100 185.000 92.500 ;
        RECT 185.400 92.400 185.800 92.800 ;
        RECT 186.300 92.700 186.700 92.800 ;
        RECT 186.300 92.400 187.700 92.700 ;
        RECT 187.400 92.100 187.700 92.400 ;
        RECT 189.400 92.100 189.800 92.500 ;
        RECT 184.600 91.800 185.600 92.100 ;
        RECT 185.200 91.100 185.600 91.800 ;
        RECT 187.400 91.100 187.800 92.100 ;
        RECT 189.400 91.800 190.100 92.100 ;
        RECT 189.500 91.100 190.100 91.800 ;
        RECT 191.800 91.100 192.200 93.300 ;
        RECT 192.600 93.400 193.700 93.700 ;
        RECT 192.600 91.100 193.000 93.400 ;
        RECT 1.900 89.200 2.300 89.900 ;
        RECT 1.400 88.800 2.300 89.200 ;
        RECT 1.900 88.200 2.300 88.800 ;
        RECT 1.400 87.900 2.300 88.200 ;
        RECT 4.900 88.000 5.300 89.500 ;
        RECT 7.000 88.500 7.400 89.500 ;
        RECT 0.600 86.800 1.000 87.600 ;
        RECT 1.400 81.100 1.800 87.900 ;
        RECT 4.500 87.700 5.300 88.000 ;
        RECT 4.500 87.500 4.900 87.700 ;
        RECT 4.500 87.200 4.800 87.500 ;
        RECT 7.100 87.400 7.400 88.500 ;
        RECT 3.800 86.800 4.800 87.200 ;
        RECT 5.300 87.100 7.400 87.400 ;
        RECT 7.800 88.500 8.200 89.500 ;
        RECT 7.800 87.400 8.100 88.500 ;
        RECT 9.900 88.000 10.300 89.500 ;
        RECT 9.900 87.700 10.700 88.000 ;
        RECT 10.300 87.500 10.700 87.700 ;
        RECT 7.800 87.100 9.900 87.400 ;
        RECT 5.300 86.900 5.800 87.100 ;
        RECT 3.800 85.400 4.200 86.200 ;
        RECT 2.200 84.400 2.600 85.200 ;
        RECT 4.500 84.900 4.800 86.800 ;
        RECT 5.100 86.500 5.800 86.900 ;
        RECT 9.400 86.900 9.900 87.100 ;
        RECT 10.400 87.200 10.700 87.500 ;
        RECT 12.600 87.700 13.000 89.900 ;
        RECT 14.700 89.200 15.300 89.900 ;
        RECT 14.700 88.900 15.400 89.200 ;
        RECT 17.000 88.900 17.400 89.900 ;
        RECT 19.200 89.200 19.600 89.900 ;
        RECT 19.200 88.900 20.200 89.200 ;
        RECT 15.000 88.500 15.400 88.900 ;
        RECT 17.100 88.600 17.400 88.900 ;
        RECT 17.100 88.300 18.500 88.600 ;
        RECT 18.100 88.200 18.500 88.300 ;
        RECT 19.000 88.200 19.400 88.600 ;
        RECT 19.800 88.500 20.200 88.900 ;
        RECT 14.100 87.700 14.500 87.800 ;
        RECT 12.600 87.400 14.500 87.700 ;
        RECT 5.500 85.500 5.800 86.500 ;
        RECT 6.200 85.800 6.600 86.600 ;
        RECT 7.000 86.100 7.400 86.600 ;
        RECT 7.800 86.100 8.200 86.600 ;
        RECT 7.000 85.800 8.200 86.100 ;
        RECT 8.600 85.800 9.000 86.600 ;
        RECT 9.400 86.500 10.100 86.900 ;
        RECT 10.400 86.800 11.400 87.200 ;
        RECT 9.400 85.500 9.700 86.500 ;
        RECT 5.500 85.200 7.400 85.500 ;
        RECT 4.500 84.600 5.300 84.900 ;
        RECT 4.900 82.200 5.300 84.600 ;
        RECT 7.100 83.500 7.400 85.200 ;
        RECT 4.900 81.800 5.800 82.200 ;
        RECT 4.900 81.100 5.300 81.800 ;
        RECT 7.000 81.500 7.400 83.500 ;
        RECT 7.800 85.200 9.700 85.500 ;
        RECT 7.800 83.500 8.100 85.200 ;
        RECT 10.400 84.900 10.700 86.800 ;
        RECT 11.000 86.100 11.400 86.200 ;
        RECT 11.800 86.100 12.200 86.200 ;
        RECT 11.000 85.800 12.200 86.100 ;
        RECT 11.000 85.400 11.400 85.800 ;
        RECT 12.600 85.700 13.000 87.400 ;
        RECT 16.100 87.100 16.500 87.200 ;
        RECT 18.200 87.100 18.600 87.200 ;
        RECT 19.000 87.100 19.300 88.200 ;
        RECT 21.400 87.500 21.800 89.900 ;
        RECT 23.000 88.200 23.400 89.900 ;
        RECT 22.900 87.900 23.400 88.200 ;
        RECT 22.900 87.200 23.200 87.900 ;
        RECT 24.600 87.600 25.000 89.900 ;
        RECT 23.700 87.300 25.000 87.600 ;
        RECT 25.400 87.600 25.800 89.900 ;
        RECT 27.000 88.200 27.400 89.900 ;
        RECT 27.000 87.900 27.500 88.200 ;
        RECT 25.400 87.300 26.700 87.600 ;
        RECT 20.600 87.100 21.400 87.200 ;
        RECT 15.900 86.800 21.400 87.100 ;
        RECT 22.900 86.800 23.400 87.200 ;
        RECT 15.000 86.400 15.400 86.500 ;
        RECT 13.500 86.100 15.400 86.400 ;
        RECT 13.500 86.000 13.900 86.100 ;
        RECT 14.300 85.700 14.700 85.800 ;
        RECT 12.600 85.400 14.700 85.700 ;
        RECT 9.900 84.600 10.700 84.900 ;
        RECT 7.800 81.500 8.200 83.500 ;
        RECT 9.900 82.200 10.300 84.600 ;
        RECT 9.900 81.800 10.600 82.200 ;
        RECT 9.900 81.100 10.300 81.800 ;
        RECT 12.600 81.100 13.000 85.400 ;
        RECT 15.900 85.200 16.200 86.800 ;
        RECT 19.500 86.700 19.900 86.800 ;
        RECT 19.000 86.200 19.400 86.300 ;
        RECT 20.300 86.200 20.700 86.300 ;
        RECT 18.200 85.900 20.700 86.200 ;
        RECT 18.200 85.800 18.600 85.900 ;
        RECT 19.000 85.500 21.800 85.600 ;
        RECT 18.900 85.400 21.800 85.500 ;
        RECT 15.000 84.900 16.200 85.200 ;
        RECT 16.900 85.300 21.800 85.400 ;
        RECT 16.900 85.100 19.300 85.300 ;
        RECT 15.000 84.400 15.300 84.900 ;
        RECT 14.600 84.000 15.300 84.400 ;
        RECT 16.100 84.500 16.500 84.600 ;
        RECT 16.900 84.500 17.200 85.100 ;
        RECT 16.100 84.200 17.200 84.500 ;
        RECT 17.500 84.500 20.200 84.800 ;
        RECT 17.500 84.400 17.900 84.500 ;
        RECT 19.800 84.400 20.200 84.500 ;
        RECT 16.700 83.700 17.100 83.800 ;
        RECT 18.100 83.700 18.500 83.800 ;
        RECT 15.000 83.100 15.400 83.500 ;
        RECT 16.700 83.400 18.500 83.700 ;
        RECT 17.100 83.100 17.400 83.400 ;
        RECT 19.800 83.100 20.200 83.500 ;
        RECT 14.700 81.100 15.300 83.100 ;
        RECT 17.000 81.100 17.400 83.100 ;
        RECT 19.200 82.800 20.200 83.100 ;
        RECT 19.200 81.100 19.600 82.800 ;
        RECT 21.400 81.100 21.800 85.300 ;
        RECT 22.900 85.100 23.200 86.800 ;
        RECT 23.700 86.500 24.000 87.300 ;
        RECT 23.500 86.100 24.000 86.500 ;
        RECT 23.700 85.100 24.000 86.100 ;
        RECT 24.500 86.200 24.900 86.600 ;
        RECT 25.500 86.200 25.900 86.600 ;
        RECT 24.500 86.100 25.000 86.200 ;
        RECT 25.400 86.100 25.900 86.200 ;
        RECT 24.500 85.800 25.900 86.100 ;
        RECT 26.400 86.500 26.700 87.300 ;
        RECT 27.200 87.200 27.500 87.900 ;
        RECT 27.000 86.800 27.500 87.200 ;
        RECT 27.800 87.100 28.200 87.200 ;
        RECT 28.600 87.100 29.000 87.600 ;
        RECT 27.800 86.800 29.000 87.100 ;
        RECT 26.400 86.100 26.900 86.500 ;
        RECT 26.400 85.100 26.700 86.100 ;
        RECT 27.200 85.100 27.500 86.800 ;
        RECT 22.900 84.600 23.400 85.100 ;
        RECT 23.700 84.800 25.000 85.100 ;
        RECT 23.000 81.100 23.400 84.600 ;
        RECT 24.600 81.100 25.000 84.800 ;
        RECT 25.400 84.800 26.700 85.100 ;
        RECT 25.400 81.100 25.800 84.800 ;
        RECT 27.000 84.600 27.500 85.100 ;
        RECT 29.400 86.100 29.800 89.900 ;
        RECT 31.000 88.900 31.400 89.900 ;
        RECT 33.900 89.200 34.300 89.900 ;
        RECT 31.000 87.200 31.300 88.900 ;
        RECT 33.900 88.800 34.600 89.200 ;
        RECT 31.800 87.800 32.200 88.600 ;
        RECT 33.900 88.200 34.300 88.800 ;
        RECT 33.400 87.900 34.300 88.200 ;
        RECT 30.200 86.800 30.600 87.200 ;
        RECT 31.000 87.100 31.400 87.200 ;
        RECT 32.600 87.100 33.000 87.600 ;
        RECT 31.000 86.800 33.000 87.100 ;
        RECT 30.200 86.200 30.500 86.800 ;
        RECT 30.200 86.100 30.600 86.200 ;
        RECT 29.400 85.800 30.600 86.100 ;
        RECT 27.000 81.100 27.400 84.600 ;
        RECT 29.400 81.100 29.800 85.800 ;
        RECT 30.200 85.400 30.600 85.800 ;
        RECT 31.000 85.100 31.300 86.800 ;
        RECT 30.500 84.700 31.400 85.100 ;
        RECT 30.500 81.100 30.900 84.700 ;
        RECT 33.400 81.100 33.800 87.900 ;
        RECT 35.000 87.800 35.400 88.600 ;
        RECT 35.000 87.200 35.300 87.800 ;
        RECT 35.000 86.800 35.400 87.200 ;
        RECT 34.200 84.400 34.600 85.200 ;
        RECT 35.000 85.100 35.400 85.200 ;
        RECT 35.800 85.100 36.200 89.900 ;
        RECT 37.900 88.200 38.300 89.900 ;
        RECT 40.300 89.200 40.700 89.900 ;
        RECT 39.800 88.800 40.700 89.200 ;
        RECT 40.300 88.200 40.700 88.800 ;
        RECT 37.400 87.800 38.500 88.200 ;
        RECT 36.600 86.800 37.000 87.600 ;
        RECT 35.000 84.800 36.200 85.100 ;
        RECT 35.800 81.100 36.200 84.800 ;
        RECT 37.400 81.100 37.800 87.800 ;
        RECT 38.200 87.200 38.500 87.800 ;
        RECT 39.800 87.900 40.700 88.200 ;
        RECT 41.400 87.900 41.800 89.900 ;
        RECT 42.200 88.000 42.600 89.900 ;
        RECT 43.800 88.000 44.200 89.900 ;
        RECT 45.400 88.800 45.800 89.900 ;
        RECT 42.200 87.900 44.200 88.000 ;
        RECT 38.200 86.800 38.600 87.200 ;
        RECT 39.000 86.800 39.400 87.600 ;
        RECT 38.200 84.400 38.600 85.200 ;
        RECT 39.800 81.100 40.200 87.900 ;
        RECT 41.500 87.200 41.800 87.900 ;
        RECT 42.300 87.700 44.100 87.900 ;
        RECT 44.600 87.800 45.000 88.600 ;
        RECT 43.400 87.200 43.800 87.400 ;
        RECT 45.500 87.200 45.800 88.800 ;
        RECT 48.600 87.900 49.000 89.900 ;
        RECT 50.800 89.200 51.600 89.900 ;
        RECT 50.800 88.800 52.200 89.200 ;
        RECT 50.800 88.100 51.600 88.800 ;
        RECT 48.600 87.600 49.900 87.900 ;
        RECT 49.500 87.500 49.900 87.600 ;
        RECT 50.200 87.400 51.000 87.800 ;
        RECT 41.400 86.800 42.700 87.200 ;
        RECT 43.400 86.900 44.200 87.200 ;
        RECT 43.800 86.800 44.200 86.900 ;
        RECT 45.400 86.800 45.800 87.200 ;
        RECT 48.600 87.100 49.400 87.200 ;
        RECT 51.300 87.100 51.600 88.100 ;
        RECT 53.400 87.900 53.800 89.900 ;
        RECT 54.200 87.900 54.600 89.900 ;
        RECT 55.000 88.000 55.400 89.900 ;
        RECT 56.600 88.000 57.000 89.900 ;
        RECT 55.000 87.900 57.000 88.000 ;
        RECT 51.900 87.400 52.300 87.800 ;
        RECT 52.600 87.600 53.800 87.900 ;
        RECT 52.600 87.500 53.000 87.600 ;
        RECT 48.600 87.000 49.700 87.100 ;
        RECT 48.600 86.800 50.800 87.000 ;
        RECT 40.600 84.400 41.000 85.200 ;
        RECT 41.400 85.100 41.800 85.200 ;
        RECT 42.400 85.100 42.700 86.800 ;
        RECT 43.000 85.800 43.400 86.600 ;
        RECT 45.500 85.100 45.800 86.800 ;
        RECT 49.400 86.700 50.800 86.800 ;
        RECT 50.400 86.600 50.800 86.700 ;
        RECT 51.100 86.800 51.600 87.100 ;
        RECT 52.000 87.200 52.300 87.400 ;
        RECT 54.300 87.200 54.600 87.900 ;
        RECT 55.100 87.700 56.900 87.900 ;
        RECT 56.200 87.200 56.600 87.400 ;
        RECT 52.000 86.800 52.400 87.200 ;
        RECT 53.000 86.800 53.800 87.200 ;
        RECT 54.200 86.800 55.500 87.200 ;
        RECT 56.200 87.100 57.000 87.200 ;
        RECT 57.400 87.100 57.800 89.900 ;
        RECT 58.200 87.800 58.600 88.600 ;
        RECT 56.200 86.900 57.800 87.100 ;
        RECT 60.800 87.100 61.200 89.900 ;
        RECT 62.200 87.700 62.600 89.900 ;
        RECT 64.300 89.200 64.900 89.900 ;
        RECT 64.300 88.900 65.000 89.200 ;
        RECT 66.600 88.900 67.000 89.900 ;
        RECT 68.800 89.200 69.200 89.900 ;
        RECT 68.800 88.900 69.800 89.200 ;
        RECT 64.600 88.500 65.000 88.900 ;
        RECT 66.700 88.600 67.000 88.900 ;
        RECT 66.700 88.300 68.100 88.600 ;
        RECT 67.700 88.200 68.100 88.300 ;
        RECT 68.600 88.200 69.000 88.600 ;
        RECT 69.400 88.500 69.800 88.900 ;
        RECT 63.700 87.700 64.100 87.800 ;
        RECT 62.200 87.400 64.100 87.700 ;
        RECT 60.800 86.900 61.700 87.100 ;
        RECT 56.600 86.800 57.800 86.900 ;
        RECT 60.900 86.800 61.700 86.900 ;
        RECT 51.100 86.200 51.400 86.800 ;
        RECT 46.200 85.400 46.600 86.200 ;
        RECT 49.700 86.100 50.100 86.200 ;
        RECT 49.700 85.800 50.500 86.100 ;
        RECT 51.000 85.800 51.400 86.200 ;
        RECT 50.100 85.700 50.500 85.800 ;
        RECT 51.100 85.100 51.400 85.800 ;
        RECT 54.200 85.100 54.600 85.200 ;
        RECT 55.200 85.100 55.500 86.800 ;
        RECT 55.800 86.100 56.200 86.600 ;
        RECT 56.600 86.100 57.000 86.200 ;
        RECT 55.800 85.800 57.000 86.100 ;
        RECT 41.400 84.800 42.100 85.100 ;
        RECT 42.400 84.800 42.900 85.100 ;
        RECT 41.800 84.200 42.100 84.800 ;
        RECT 42.500 84.200 42.900 84.800 ;
        RECT 45.400 84.700 46.300 85.100 ;
        RECT 41.800 83.800 42.200 84.200 ;
        RECT 42.500 83.800 43.400 84.200 ;
        RECT 42.500 81.100 42.900 83.800 ;
        RECT 45.900 81.100 46.300 84.700 ;
        RECT 48.600 84.800 49.900 85.100 ;
        RECT 48.600 81.100 49.000 84.800 ;
        RECT 49.500 84.700 49.900 84.800 ;
        RECT 50.800 81.100 51.600 85.100 ;
        RECT 52.600 84.800 53.800 85.100 ;
        RECT 54.200 84.800 54.900 85.100 ;
        RECT 55.200 84.800 55.700 85.100 ;
        RECT 52.600 84.700 53.000 84.800 ;
        RECT 53.400 81.100 53.800 84.800 ;
        RECT 54.600 84.200 54.900 84.800 ;
        RECT 54.600 83.800 55.000 84.200 ;
        RECT 55.300 81.100 55.700 84.800 ;
        RECT 57.400 81.100 57.800 86.800 ;
        RECT 59.800 85.800 60.600 86.200 ;
        RECT 59.000 84.800 59.400 85.600 ;
        RECT 61.400 85.200 61.700 86.800 ;
        RECT 62.200 85.700 62.600 87.400 ;
        RECT 65.700 87.100 66.100 87.200 ;
        RECT 68.600 87.100 68.900 88.200 ;
        RECT 71.000 87.500 71.400 89.900 ;
        RECT 72.100 89.200 72.500 89.900 ;
        RECT 72.100 88.800 73.000 89.200 ;
        RECT 72.100 88.200 72.500 88.800 ;
        RECT 72.100 87.900 73.000 88.200 ;
        RECT 70.200 87.100 71.000 87.200 ;
        RECT 65.500 86.800 71.000 87.100 ;
        RECT 64.600 86.400 65.000 86.500 ;
        RECT 63.100 86.100 65.000 86.400 ;
        RECT 63.100 86.000 63.500 86.100 ;
        RECT 63.900 85.700 64.300 85.800 ;
        RECT 62.200 85.400 64.300 85.700 ;
        RECT 61.400 84.800 61.800 85.200 ;
        RECT 59.800 84.100 60.200 84.200 ;
        RECT 60.600 84.100 61.000 84.600 ;
        RECT 59.800 83.800 61.000 84.100 ;
        RECT 61.400 83.500 61.700 84.800 ;
        RECT 59.900 83.200 61.700 83.500 ;
        RECT 59.900 83.100 60.200 83.200 ;
        RECT 59.800 81.100 60.200 83.100 ;
        RECT 61.400 83.100 61.700 83.200 ;
        RECT 61.400 81.100 61.800 83.100 ;
        RECT 62.200 81.100 62.600 85.400 ;
        RECT 65.500 85.200 65.800 86.800 ;
        RECT 69.100 86.700 69.500 86.800 ;
        RECT 68.600 86.200 69.000 86.300 ;
        RECT 69.900 86.200 70.300 86.300 ;
        RECT 67.800 85.900 70.300 86.200 ;
        RECT 67.800 85.800 68.200 85.900 ;
        RECT 68.600 85.500 71.400 85.600 ;
        RECT 68.500 85.400 71.400 85.500 ;
        RECT 64.600 84.900 65.800 85.200 ;
        RECT 66.500 85.300 71.400 85.400 ;
        RECT 66.500 85.100 68.900 85.300 ;
        RECT 64.600 84.400 64.900 84.900 ;
        RECT 64.200 84.000 64.900 84.400 ;
        RECT 65.700 84.500 66.100 84.600 ;
        RECT 66.500 84.500 66.800 85.100 ;
        RECT 65.700 84.200 66.800 84.500 ;
        RECT 67.100 84.500 69.800 84.800 ;
        RECT 67.100 84.400 67.500 84.500 ;
        RECT 69.400 84.400 69.800 84.500 ;
        RECT 66.300 83.700 66.700 83.800 ;
        RECT 67.700 83.700 68.100 83.800 ;
        RECT 64.600 83.100 65.000 83.500 ;
        RECT 66.300 83.400 68.100 83.700 ;
        RECT 66.700 83.100 67.000 83.400 ;
        RECT 69.400 83.100 69.800 83.500 ;
        RECT 64.300 81.100 64.900 83.100 ;
        RECT 66.600 81.100 67.000 83.100 ;
        RECT 68.800 82.800 69.800 83.100 ;
        RECT 68.800 81.100 69.200 82.800 ;
        RECT 71.000 81.100 71.400 85.300 ;
        RECT 71.800 84.400 72.200 85.200 ;
        RECT 72.600 81.100 73.000 87.900 ;
        RECT 74.200 87.700 74.600 89.900 ;
        RECT 76.300 89.200 76.900 89.900 ;
        RECT 76.300 88.900 77.000 89.200 ;
        RECT 78.600 88.900 79.000 89.900 ;
        RECT 80.800 89.200 81.200 89.900 ;
        RECT 80.800 88.900 81.800 89.200 ;
        RECT 76.600 88.500 77.000 88.900 ;
        RECT 78.700 88.600 79.000 88.900 ;
        RECT 78.700 88.300 80.100 88.600 ;
        RECT 79.700 88.200 80.100 88.300 ;
        RECT 80.600 88.200 81.000 88.600 ;
        RECT 81.400 88.500 81.800 88.900 ;
        RECT 75.700 87.700 76.100 87.800 ;
        RECT 73.400 87.100 73.800 87.600 ;
        RECT 74.200 87.400 76.100 87.700 ;
        RECT 74.200 87.100 74.600 87.400 ;
        RECT 77.700 87.100 78.100 87.200 ;
        RECT 80.600 87.100 80.900 88.200 ;
        RECT 83.000 87.500 83.400 89.900 ;
        RECT 84.600 88.200 85.000 89.900 ;
        RECT 84.500 87.900 85.000 88.200 ;
        RECT 84.500 87.200 84.800 87.900 ;
        RECT 86.200 87.600 86.600 89.900 ;
        RECT 85.300 87.300 86.600 87.600 ;
        RECT 87.000 87.700 87.400 89.900 ;
        RECT 89.100 89.200 89.700 89.900 ;
        RECT 89.100 88.900 89.800 89.200 ;
        RECT 91.400 88.900 91.800 89.900 ;
        RECT 93.600 89.200 94.000 89.900 ;
        RECT 93.600 88.900 94.600 89.200 ;
        RECT 89.400 88.500 89.800 88.900 ;
        RECT 91.500 88.600 91.800 88.900 ;
        RECT 91.500 88.300 92.900 88.600 ;
        RECT 92.500 88.200 92.900 88.300 ;
        RECT 93.400 88.200 93.800 88.600 ;
        RECT 94.200 88.500 94.600 88.900 ;
        RECT 88.500 87.700 88.900 87.800 ;
        RECT 87.000 87.400 88.900 87.700 ;
        RECT 82.200 87.100 83.000 87.200 ;
        RECT 73.400 86.800 74.600 87.100 ;
        RECT 74.200 85.700 74.600 86.800 ;
        RECT 77.500 86.800 83.000 87.100 ;
        RECT 84.500 86.800 85.000 87.200 ;
        RECT 76.600 86.400 77.000 86.500 ;
        RECT 75.100 86.100 77.000 86.400 ;
        RECT 75.100 86.000 75.500 86.100 ;
        RECT 75.900 85.700 76.300 85.800 ;
        RECT 74.200 85.400 76.300 85.700 ;
        RECT 74.200 81.100 74.600 85.400 ;
        RECT 77.500 85.200 77.800 86.800 ;
        RECT 81.100 86.700 81.500 86.800 ;
        RECT 81.900 86.200 82.300 86.300 ;
        RECT 79.000 86.100 79.400 86.200 ;
        RECT 79.800 86.100 82.300 86.200 ;
        RECT 79.000 85.900 82.300 86.100 ;
        RECT 79.000 85.800 80.200 85.900 ;
        RECT 80.600 85.500 83.400 85.600 ;
        RECT 80.500 85.400 83.400 85.500 ;
        RECT 76.600 84.900 77.800 85.200 ;
        RECT 78.500 85.300 83.400 85.400 ;
        RECT 78.500 85.100 80.900 85.300 ;
        RECT 76.600 84.400 76.900 84.900 ;
        RECT 76.200 84.000 76.900 84.400 ;
        RECT 77.700 84.500 78.100 84.600 ;
        RECT 78.500 84.500 78.800 85.100 ;
        RECT 77.700 84.200 78.800 84.500 ;
        RECT 79.100 84.500 81.800 84.800 ;
        RECT 79.100 84.400 79.500 84.500 ;
        RECT 81.400 84.400 81.800 84.500 ;
        RECT 78.300 83.700 78.700 83.800 ;
        RECT 79.700 83.700 80.100 83.800 ;
        RECT 76.600 83.100 77.000 83.500 ;
        RECT 78.300 83.400 80.100 83.700 ;
        RECT 78.700 83.100 79.000 83.400 ;
        RECT 81.400 83.100 81.800 83.500 ;
        RECT 76.300 81.100 76.900 83.100 ;
        RECT 78.600 81.100 79.000 83.100 ;
        RECT 80.800 82.800 81.800 83.100 ;
        RECT 80.800 81.100 81.200 82.800 ;
        RECT 83.000 81.100 83.400 85.300 ;
        RECT 84.500 85.100 84.800 86.800 ;
        RECT 85.300 86.500 85.600 87.300 ;
        RECT 85.100 86.100 85.600 86.500 ;
        RECT 85.300 85.100 85.600 86.100 ;
        RECT 86.100 86.200 86.500 86.600 ;
        RECT 86.100 85.800 86.600 86.200 ;
        RECT 87.000 85.700 87.400 87.400 ;
        RECT 90.500 87.100 90.900 87.200 ;
        RECT 93.400 87.100 93.700 88.200 ;
        RECT 95.800 87.500 96.200 89.900 ;
        RECT 98.200 87.700 98.600 89.900 ;
        RECT 100.300 89.200 100.900 89.900 ;
        RECT 100.300 88.900 101.000 89.200 ;
        RECT 102.600 88.900 103.000 89.900 ;
        RECT 104.800 89.200 105.200 89.900 ;
        RECT 104.800 88.900 105.800 89.200 ;
        RECT 100.600 88.500 101.000 88.900 ;
        RECT 102.700 88.600 103.000 88.900 ;
        RECT 102.700 88.300 104.100 88.600 ;
        RECT 103.700 88.200 104.100 88.300 ;
        RECT 104.600 88.200 105.000 88.600 ;
        RECT 105.400 88.500 105.800 88.900 ;
        RECT 99.700 87.700 100.100 87.800 ;
        RECT 98.200 87.400 100.100 87.700 ;
        RECT 95.000 87.100 95.800 87.200 ;
        RECT 90.300 86.800 95.800 87.100 ;
        RECT 89.400 86.400 89.800 86.500 ;
        RECT 87.900 86.100 89.800 86.400 ;
        RECT 87.900 86.000 88.300 86.100 ;
        RECT 88.700 85.700 89.100 85.800 ;
        RECT 87.000 85.400 89.100 85.700 ;
        RECT 84.500 84.600 85.000 85.100 ;
        RECT 85.300 84.800 86.600 85.100 ;
        RECT 84.600 81.100 85.000 84.600 ;
        RECT 86.200 81.100 86.600 84.800 ;
        RECT 87.000 81.100 87.400 85.400 ;
        RECT 90.300 85.200 90.600 86.800 ;
        RECT 93.900 86.700 94.300 86.800 ;
        RECT 93.400 86.200 93.800 86.300 ;
        RECT 94.700 86.200 95.100 86.300 ;
        RECT 92.600 85.900 95.100 86.200 ;
        RECT 92.600 85.800 93.000 85.900 ;
        RECT 98.200 85.700 98.600 87.400 ;
        RECT 101.700 87.100 102.100 87.200 ;
        RECT 104.600 87.100 104.900 88.200 ;
        RECT 107.000 87.500 107.400 89.900 ;
        RECT 107.800 87.700 108.200 89.900 ;
        RECT 109.900 89.200 110.500 89.900 ;
        RECT 109.900 88.900 110.600 89.200 ;
        RECT 112.200 88.900 112.600 89.900 ;
        RECT 114.400 89.200 114.800 89.900 ;
        RECT 114.400 88.900 115.400 89.200 ;
        RECT 110.200 88.500 110.600 88.900 ;
        RECT 112.300 88.600 112.600 88.900 ;
        RECT 112.300 88.300 113.700 88.600 ;
        RECT 113.300 88.200 113.700 88.300 ;
        RECT 114.200 88.200 114.600 88.600 ;
        RECT 115.000 88.500 115.400 88.900 ;
        RECT 109.400 87.800 109.800 88.200 ;
        RECT 109.300 87.700 109.800 87.800 ;
        RECT 107.800 87.400 109.800 87.700 ;
        RECT 106.200 87.100 107.000 87.200 ;
        RECT 101.500 86.800 107.000 87.100 ;
        RECT 100.600 86.400 101.000 86.500 ;
        RECT 99.100 86.100 101.000 86.400 ;
        RECT 99.100 86.000 99.500 86.100 ;
        RECT 99.900 85.700 100.300 85.800 ;
        RECT 93.400 85.500 96.200 85.600 ;
        RECT 93.300 85.400 96.200 85.500 ;
        RECT 89.400 84.900 90.600 85.200 ;
        RECT 91.300 85.300 96.200 85.400 ;
        RECT 91.300 85.100 93.700 85.300 ;
        RECT 89.400 84.400 89.700 84.900 ;
        RECT 89.000 84.200 89.700 84.400 ;
        RECT 90.500 84.500 90.900 84.600 ;
        RECT 91.300 84.500 91.600 85.100 ;
        RECT 90.500 84.200 91.600 84.500 ;
        RECT 91.900 84.500 94.600 84.800 ;
        RECT 91.900 84.400 92.300 84.500 ;
        RECT 94.200 84.400 94.600 84.500 ;
        RECT 88.600 84.000 89.700 84.200 ;
        RECT 88.600 83.800 89.300 84.000 ;
        RECT 91.100 83.700 91.500 83.800 ;
        RECT 92.500 83.700 92.900 83.800 ;
        RECT 89.400 83.100 89.800 83.500 ;
        RECT 91.100 83.400 92.900 83.700 ;
        RECT 91.500 83.100 91.800 83.400 ;
        RECT 94.200 83.100 94.600 83.500 ;
        RECT 89.100 81.100 89.700 83.100 ;
        RECT 91.400 81.100 91.800 83.100 ;
        RECT 93.600 82.800 94.600 83.100 ;
        RECT 93.600 81.100 94.000 82.800 ;
        RECT 95.800 81.100 96.200 85.300 ;
        RECT 98.200 85.400 100.300 85.700 ;
        RECT 98.200 81.100 98.600 85.400 ;
        RECT 101.500 85.200 101.800 86.800 ;
        RECT 105.100 86.700 105.500 86.800 ;
        RECT 104.600 86.200 105.000 86.300 ;
        RECT 105.900 86.200 106.300 86.300 ;
        RECT 103.800 85.900 106.300 86.200 ;
        RECT 103.800 85.800 104.200 85.900 ;
        RECT 107.800 85.700 108.200 87.400 ;
        RECT 111.300 87.100 111.700 87.200 ;
        RECT 114.200 87.100 114.500 88.200 ;
        RECT 116.600 87.500 117.000 89.900 ;
        RECT 118.200 88.900 118.600 89.900 ;
        RECT 117.400 87.800 117.800 88.600 ;
        RECT 118.300 87.200 118.600 88.900 ;
        RECT 120.100 89.200 120.500 89.900 ;
        RECT 120.100 88.800 121.000 89.200 ;
        RECT 120.100 88.200 120.500 88.800 ;
        RECT 122.200 88.500 122.600 89.500 ;
        RECT 120.100 87.900 121.000 88.200 ;
        RECT 115.800 87.100 116.600 87.200 ;
        RECT 111.100 86.800 116.600 87.100 ;
        RECT 118.200 86.800 118.600 87.200 ;
        RECT 110.200 86.400 110.600 86.500 ;
        RECT 108.700 86.100 110.600 86.400 ;
        RECT 111.100 86.200 111.400 86.800 ;
        RECT 114.700 86.700 115.100 86.800 ;
        RECT 115.500 86.200 115.900 86.300 ;
        RECT 108.700 86.000 109.100 86.100 ;
        RECT 111.000 85.800 111.400 86.200 ;
        RECT 113.400 85.900 115.900 86.200 ;
        RECT 113.400 85.800 113.800 85.900 ;
        RECT 109.500 85.700 109.900 85.800 ;
        RECT 104.600 85.500 107.400 85.600 ;
        RECT 104.500 85.400 107.400 85.500 ;
        RECT 100.600 84.900 101.800 85.200 ;
        RECT 102.500 85.300 107.400 85.400 ;
        RECT 102.500 85.100 104.900 85.300 ;
        RECT 100.600 84.400 100.900 84.900 ;
        RECT 100.200 84.000 100.900 84.400 ;
        RECT 101.700 84.500 102.100 84.600 ;
        RECT 102.500 84.500 102.800 85.100 ;
        RECT 101.700 84.200 102.800 84.500 ;
        RECT 103.100 84.500 105.800 84.800 ;
        RECT 103.100 84.400 103.500 84.500 ;
        RECT 105.400 84.400 105.800 84.500 ;
        RECT 102.300 83.700 102.700 83.800 ;
        RECT 103.700 83.700 104.100 83.800 ;
        RECT 100.600 83.100 101.000 83.500 ;
        RECT 102.300 83.400 104.100 83.700 ;
        RECT 102.700 83.100 103.000 83.400 ;
        RECT 105.400 83.100 105.800 83.500 ;
        RECT 100.300 81.100 100.900 83.100 ;
        RECT 102.600 81.100 103.000 83.100 ;
        RECT 104.800 82.800 105.800 83.100 ;
        RECT 104.800 81.100 105.200 82.800 ;
        RECT 107.000 81.100 107.400 85.300 ;
        RECT 107.800 85.400 109.900 85.700 ;
        RECT 107.800 81.100 108.200 85.400 ;
        RECT 111.100 85.200 111.400 85.800 ;
        RECT 114.200 85.500 117.000 85.600 ;
        RECT 114.100 85.400 117.000 85.500 ;
        RECT 110.200 84.900 111.400 85.200 ;
        RECT 112.100 85.300 117.000 85.400 ;
        RECT 112.100 85.100 114.500 85.300 ;
        RECT 110.200 84.400 110.500 84.900 ;
        RECT 109.800 84.000 110.500 84.400 ;
        RECT 111.300 84.500 111.700 84.600 ;
        RECT 112.100 84.500 112.400 85.100 ;
        RECT 111.300 84.200 112.400 84.500 ;
        RECT 112.700 84.500 115.400 84.800 ;
        RECT 112.700 84.400 113.100 84.500 ;
        RECT 115.000 84.400 115.400 84.500 ;
        RECT 111.900 83.700 112.300 83.800 ;
        RECT 113.300 83.700 113.700 83.800 ;
        RECT 110.200 83.100 110.600 83.500 ;
        RECT 111.900 83.400 113.700 83.700 ;
        RECT 112.300 83.100 112.600 83.400 ;
        RECT 115.000 83.100 115.400 83.500 ;
        RECT 109.900 81.100 110.500 83.100 ;
        RECT 112.200 81.100 112.600 83.100 ;
        RECT 114.400 82.800 115.400 83.100 ;
        RECT 114.400 81.100 114.800 82.800 ;
        RECT 116.600 81.100 117.000 85.300 ;
        RECT 118.300 85.100 118.600 86.800 ;
        RECT 119.000 85.400 119.400 86.200 ;
        RECT 118.200 84.700 119.100 85.100 ;
        RECT 118.700 82.200 119.100 84.700 ;
        RECT 119.800 84.400 120.200 85.200 ;
        RECT 118.700 81.800 119.400 82.200 ;
        RECT 118.700 81.100 119.100 81.800 ;
        RECT 120.600 81.100 121.000 87.900 ;
        RECT 121.400 86.800 121.800 87.600 ;
        RECT 122.200 87.400 122.500 88.500 ;
        RECT 124.300 88.200 124.700 89.500 ;
        RECT 123.800 88.000 124.700 88.200 ;
        RECT 123.800 87.800 125.100 88.000 ;
        RECT 124.300 87.700 125.100 87.800 ;
        RECT 124.700 87.500 125.100 87.700 ;
        RECT 122.200 87.100 124.300 87.400 ;
        RECT 123.800 86.900 124.300 87.100 ;
        RECT 124.800 87.200 125.100 87.500 ;
        RECT 127.000 87.700 127.400 89.900 ;
        RECT 129.100 89.200 129.700 89.900 ;
        RECT 129.100 88.900 129.800 89.200 ;
        RECT 131.400 88.900 131.800 89.900 ;
        RECT 133.600 89.200 134.000 89.900 ;
        RECT 133.600 88.900 134.600 89.200 ;
        RECT 129.400 88.500 129.800 88.900 ;
        RECT 131.500 88.600 131.800 88.900 ;
        RECT 131.500 88.300 132.900 88.600 ;
        RECT 132.500 88.200 132.900 88.300 ;
        RECT 133.400 88.200 133.800 88.600 ;
        RECT 134.200 88.500 134.600 88.900 ;
        RECT 128.500 87.700 128.900 87.800 ;
        RECT 127.000 87.400 128.900 87.700 ;
        RECT 122.200 85.800 122.600 86.600 ;
        RECT 123.000 85.800 123.400 86.600 ;
        RECT 123.800 86.500 124.500 86.900 ;
        RECT 124.800 86.800 125.800 87.200 ;
        RECT 123.800 85.500 124.100 86.500 ;
        RECT 122.200 85.200 124.100 85.500 ;
        RECT 122.200 83.500 122.500 85.200 ;
        RECT 124.800 84.900 125.100 86.800 ;
        RECT 125.400 85.400 125.800 86.200 ;
        RECT 127.000 85.700 127.400 87.400 ;
        RECT 133.400 87.200 133.700 88.200 ;
        RECT 135.800 87.500 136.200 89.900 ;
        RECT 137.400 88.900 137.800 89.900 ;
        RECT 136.600 87.800 137.000 88.600 ;
        RECT 137.500 87.200 137.800 88.900 ;
        RECT 140.900 88.000 141.300 89.500 ;
        RECT 143.000 88.500 143.400 89.500 ;
        RECT 140.500 87.700 141.300 88.000 ;
        RECT 140.500 87.500 140.900 87.700 ;
        RECT 140.500 87.200 140.800 87.500 ;
        RECT 143.100 87.400 143.400 88.500 ;
        RECT 130.500 87.100 130.900 87.200 ;
        RECT 133.400 87.100 133.800 87.200 ;
        RECT 135.000 87.100 135.800 87.200 ;
        RECT 130.300 86.800 135.800 87.100 ;
        RECT 137.400 87.100 137.800 87.200 ;
        RECT 138.200 87.100 138.600 87.200 ;
        RECT 137.400 86.800 138.600 87.100 ;
        RECT 139.000 86.800 139.400 87.200 ;
        RECT 139.800 86.800 140.800 87.200 ;
        RECT 141.300 87.100 143.400 87.400 ;
        RECT 145.400 87.700 145.800 89.900 ;
        RECT 147.500 89.200 148.100 89.900 ;
        RECT 147.500 88.900 148.200 89.200 ;
        RECT 149.800 88.900 150.200 89.900 ;
        RECT 152.000 89.200 152.400 89.900 ;
        RECT 152.000 88.900 153.000 89.200 ;
        RECT 147.800 88.500 148.200 88.900 ;
        RECT 149.900 88.600 150.200 88.900 ;
        RECT 149.900 88.300 151.300 88.600 ;
        RECT 150.900 88.200 151.300 88.300 ;
        RECT 151.800 88.200 152.200 88.600 ;
        RECT 152.600 88.500 153.000 88.900 ;
        RECT 146.900 87.700 147.300 87.800 ;
        RECT 145.400 87.400 147.300 87.700 ;
        RECT 141.300 86.900 141.800 87.100 ;
        RECT 129.400 86.400 129.800 86.500 ;
        RECT 127.900 86.100 129.800 86.400 ;
        RECT 127.900 86.000 128.300 86.100 ;
        RECT 128.700 85.700 129.100 85.800 ;
        RECT 127.000 85.400 129.100 85.700 ;
        RECT 124.300 84.600 125.100 84.900 ;
        RECT 122.200 81.500 122.600 83.500 ;
        RECT 124.300 81.100 124.700 84.600 ;
        RECT 127.000 81.100 127.400 85.400 ;
        RECT 130.300 85.200 130.600 86.800 ;
        RECT 133.900 86.700 134.300 86.800 ;
        RECT 134.700 86.200 135.100 86.300 ;
        RECT 132.600 85.900 135.100 86.200 ;
        RECT 132.600 85.800 133.000 85.900 ;
        RECT 133.400 85.500 136.200 85.600 ;
        RECT 133.300 85.400 136.200 85.500 ;
        RECT 129.400 84.900 130.600 85.200 ;
        RECT 131.300 85.300 136.200 85.400 ;
        RECT 131.300 85.100 133.700 85.300 ;
        RECT 129.400 84.400 129.700 84.900 ;
        RECT 129.000 84.000 129.700 84.400 ;
        RECT 130.500 84.500 130.900 84.600 ;
        RECT 131.300 84.500 131.600 85.100 ;
        RECT 130.500 84.200 131.600 84.500 ;
        RECT 131.900 84.500 134.600 84.800 ;
        RECT 131.900 84.400 132.300 84.500 ;
        RECT 134.200 84.400 134.600 84.500 ;
        RECT 131.100 83.700 131.500 83.800 ;
        RECT 132.500 83.700 132.900 83.800 ;
        RECT 129.400 83.100 129.800 83.500 ;
        RECT 131.100 83.400 132.900 83.700 ;
        RECT 131.500 83.100 131.800 83.400 ;
        RECT 134.200 83.100 134.600 83.500 ;
        RECT 129.100 81.100 129.700 83.100 ;
        RECT 131.400 81.100 131.800 83.100 ;
        RECT 133.600 82.800 134.600 83.100 ;
        RECT 133.600 81.100 134.000 82.800 ;
        RECT 135.800 81.100 136.200 85.300 ;
        RECT 137.500 85.100 137.800 86.800 ;
        RECT 138.200 85.400 138.600 86.200 ;
        RECT 139.000 86.100 139.300 86.800 ;
        RECT 139.800 86.100 140.200 86.200 ;
        RECT 139.000 85.800 140.200 86.100 ;
        RECT 139.800 85.400 140.200 85.800 ;
        RECT 140.500 85.200 140.800 86.800 ;
        RECT 141.100 86.500 141.800 86.900 ;
        RECT 141.500 85.500 141.800 86.500 ;
        RECT 142.200 85.800 142.600 86.600 ;
        RECT 143.000 85.800 143.400 86.600 ;
        RECT 145.400 85.700 145.800 87.400 ;
        RECT 148.900 87.100 149.300 87.200 ;
        RECT 151.000 87.100 151.400 87.200 ;
        RECT 151.800 87.100 152.100 88.200 ;
        RECT 154.200 87.500 154.600 89.900 ;
        RECT 155.000 87.600 155.400 89.900 ;
        RECT 155.000 87.300 156.100 87.600 ;
        RECT 153.400 87.100 154.200 87.200 ;
        RECT 148.700 86.800 154.200 87.100 ;
        RECT 147.800 86.400 148.200 86.500 ;
        RECT 146.300 86.100 148.200 86.400 ;
        RECT 146.300 86.000 146.700 86.100 ;
        RECT 147.100 85.700 147.500 85.800 ;
        RECT 141.500 85.200 143.400 85.500 ;
        RECT 137.400 84.700 138.300 85.100 ;
        RECT 137.900 81.100 138.300 84.700 ;
        RECT 140.500 84.900 141.000 85.200 ;
        RECT 140.500 84.600 141.300 84.900 ;
        RECT 140.900 81.100 141.300 84.600 ;
        RECT 143.100 83.500 143.400 85.200 ;
        RECT 143.000 81.500 143.400 83.500 ;
        RECT 145.400 85.400 147.500 85.700 ;
        RECT 145.400 81.100 145.800 85.400 ;
        RECT 148.700 85.200 149.000 86.800 ;
        RECT 152.300 86.700 152.700 86.800 ;
        RECT 153.100 86.200 153.500 86.300 ;
        RECT 150.200 86.100 150.600 86.200 ;
        RECT 151.000 86.100 153.500 86.200 ;
        RECT 150.200 85.900 153.500 86.100 ;
        RECT 150.200 85.800 151.400 85.900 ;
        RECT 155.800 85.800 156.100 87.300 ;
        RECT 156.600 86.200 157.000 89.900 ;
        RECT 157.400 88.000 157.800 89.900 ;
        RECT 159.000 88.000 159.400 89.900 ;
        RECT 157.400 87.900 159.400 88.000 ;
        RECT 159.800 87.900 160.200 89.900 ;
        RECT 160.900 88.200 161.300 89.900 ;
        RECT 160.900 87.900 161.800 88.200 ;
        RECT 157.500 87.700 159.300 87.900 ;
        RECT 157.800 87.200 158.200 87.400 ;
        RECT 159.800 87.200 160.100 87.900 ;
        RECT 157.400 86.900 158.200 87.200 ;
        RECT 157.400 86.800 157.800 86.900 ;
        RECT 158.900 86.800 160.200 87.200 ;
        RECT 151.800 85.500 154.600 85.600 ;
        RECT 151.700 85.400 154.600 85.500 ;
        RECT 147.800 84.900 149.000 85.200 ;
        RECT 149.700 85.300 154.600 85.400 ;
        RECT 149.700 85.100 152.100 85.300 ;
        RECT 147.800 84.400 148.100 84.900 ;
        RECT 147.400 84.000 148.100 84.400 ;
        RECT 148.900 84.500 149.300 84.600 ;
        RECT 149.700 84.500 150.000 85.100 ;
        RECT 148.900 84.200 150.000 84.500 ;
        RECT 150.300 84.500 153.000 84.800 ;
        RECT 150.300 84.400 150.700 84.500 ;
        RECT 152.600 84.400 153.000 84.500 ;
        RECT 149.500 83.700 149.900 83.800 ;
        RECT 150.900 83.700 151.300 83.800 ;
        RECT 147.800 83.100 148.200 83.500 ;
        RECT 149.500 83.400 151.300 83.700 ;
        RECT 149.900 83.100 150.200 83.400 ;
        RECT 152.600 83.100 153.000 83.500 ;
        RECT 147.500 81.100 148.100 83.100 ;
        RECT 149.800 81.100 150.200 83.100 ;
        RECT 152.000 82.800 153.000 83.100 ;
        RECT 152.000 81.100 152.400 82.800 ;
        RECT 154.200 81.100 154.600 85.300 ;
        RECT 155.800 85.400 156.400 85.800 ;
        RECT 155.800 85.100 156.100 85.400 ;
        RECT 156.700 85.100 157.000 86.200 ;
        RECT 158.900 85.100 159.200 86.800 ;
        RECT 161.400 86.100 161.800 87.900 ;
        RECT 162.200 86.800 162.600 87.600 ;
        RECT 163.600 87.100 164.000 89.900 ;
        RECT 163.100 86.900 164.000 87.100 ;
        RECT 168.000 87.100 168.400 89.900 ;
        RECT 170.200 88.900 170.600 89.900 ;
        RECT 169.400 87.800 169.800 88.600 ;
        RECT 170.300 87.200 170.600 88.900 ;
        RECT 168.000 86.900 168.900 87.100 ;
        RECT 163.100 86.800 163.900 86.900 ;
        RECT 168.100 86.800 168.900 86.900 ;
        RECT 170.200 86.800 170.600 87.200 ;
        RECT 159.800 85.800 161.800 86.100 ;
        RECT 159.800 85.200 160.100 85.800 ;
        RECT 159.800 85.100 160.200 85.200 ;
        RECT 155.000 84.800 156.100 85.100 ;
        RECT 155.000 81.100 155.400 84.800 ;
        RECT 156.600 81.100 157.000 85.100 ;
        RECT 158.700 84.800 159.200 85.100 ;
        RECT 159.500 84.800 160.200 85.100 ;
        RECT 158.700 81.100 159.100 84.800 ;
        RECT 159.500 84.200 159.800 84.800 ;
        RECT 159.400 83.800 159.800 84.200 ;
        RECT 161.400 81.100 161.800 85.800 ;
        RECT 163.100 85.200 163.400 86.800 ;
        RECT 164.200 85.800 165.000 86.200 ;
        RECT 163.000 84.800 163.400 85.200 ;
        RECT 165.400 84.800 165.800 85.600 ;
        RECT 166.200 84.800 166.600 86.200 ;
        RECT 167.000 85.800 168.200 86.200 ;
        RECT 168.600 85.200 168.900 86.800 ;
        RECT 168.600 84.800 169.000 85.200 ;
        RECT 170.300 85.100 170.600 86.800 ;
        RECT 171.800 86.800 172.200 87.600 ;
        RECT 171.000 86.100 171.400 86.200 ;
        RECT 171.800 86.100 172.100 86.800 ;
        RECT 171.000 85.800 172.100 86.100 ;
        RECT 172.600 86.100 173.000 89.900 ;
        RECT 173.400 88.000 173.800 89.900 ;
        RECT 175.000 88.000 175.400 89.900 ;
        RECT 173.400 87.900 175.400 88.000 ;
        RECT 175.800 87.900 176.200 89.900 ;
        RECT 177.400 88.900 177.800 89.900 ;
        RECT 173.500 87.700 175.300 87.900 ;
        RECT 173.800 87.200 174.200 87.400 ;
        RECT 175.800 87.200 176.100 87.900 ;
        RECT 176.600 87.800 177.000 88.600 ;
        RECT 177.500 87.200 177.800 88.900 ;
        RECT 179.800 88.900 180.200 89.900 ;
        RECT 179.000 88.100 179.400 88.200 ;
        RECT 179.800 88.100 180.100 88.900 ;
        RECT 179.000 87.800 180.100 88.100 ;
        RECT 173.400 86.900 174.200 87.200 ;
        RECT 173.400 86.800 173.800 86.900 ;
        RECT 174.900 86.800 176.200 87.200 ;
        RECT 177.400 86.800 177.800 87.200 ;
        RECT 174.200 86.100 174.600 86.600 ;
        RECT 172.600 85.800 174.600 86.100 ;
        RECT 171.000 85.400 171.400 85.800 ;
        RECT 163.100 83.500 163.400 84.800 ;
        RECT 163.800 83.800 164.200 84.600 ;
        RECT 167.800 83.800 168.200 84.600 ;
        RECT 168.600 83.500 168.900 84.800 ;
        RECT 170.200 84.700 171.100 85.100 ;
        RECT 170.700 84.200 171.100 84.700 ;
        RECT 170.200 83.800 171.100 84.200 ;
        RECT 163.100 83.200 164.900 83.500 ;
        RECT 163.100 83.100 163.400 83.200 ;
        RECT 163.000 81.100 163.400 83.100 ;
        RECT 164.600 83.100 164.900 83.200 ;
        RECT 167.100 83.200 168.900 83.500 ;
        RECT 167.100 83.100 167.400 83.200 ;
        RECT 164.600 81.100 165.000 83.100 ;
        RECT 167.000 81.100 167.400 83.100 ;
        RECT 168.600 83.100 168.900 83.200 ;
        RECT 168.600 81.100 169.000 83.100 ;
        RECT 170.700 81.100 171.100 83.800 ;
        RECT 172.600 81.100 173.000 85.800 ;
        RECT 174.900 85.100 175.200 86.800 ;
        RECT 175.800 85.100 176.200 85.200 ;
        RECT 177.500 85.100 177.800 86.800 ;
        RECT 179.800 87.200 180.100 87.800 ;
        RECT 180.600 87.800 181.000 88.600 ;
        RECT 181.400 87.900 181.800 89.900 ;
        RECT 183.600 88.100 184.400 89.900 ;
        RECT 179.800 86.800 180.200 87.200 ;
        RECT 178.200 85.400 178.600 86.200 ;
        RECT 179.000 85.400 179.400 86.200 ;
        RECT 179.800 85.100 180.100 86.800 ;
        RECT 180.600 86.100 180.900 87.800 ;
        RECT 181.400 87.600 182.600 87.900 ;
        RECT 182.200 87.500 182.600 87.600 ;
        RECT 182.900 87.400 183.300 87.800 ;
        RECT 182.900 87.200 183.200 87.400 ;
        RECT 181.400 86.800 182.200 87.200 ;
        RECT 182.800 86.800 183.200 87.200 ;
        RECT 183.600 86.400 183.900 88.100 ;
        RECT 186.200 87.900 186.600 89.900 ;
        RECT 184.200 87.700 185.000 87.800 ;
        RECT 184.200 87.400 185.200 87.700 ;
        RECT 185.500 87.600 186.600 87.900 ;
        RECT 185.500 87.500 185.900 87.600 ;
        RECT 184.900 87.200 185.200 87.400 ;
        RECT 184.200 86.700 184.600 87.100 ;
        RECT 184.900 86.900 186.600 87.200 ;
        RECT 185.800 86.800 186.600 86.900 ;
        RECT 183.400 86.200 183.900 86.400 ;
        RECT 183.000 86.100 183.900 86.200 ;
        RECT 184.300 86.400 184.600 86.700 ;
        RECT 184.300 86.100 185.600 86.400 ;
        RECT 180.600 85.800 183.700 86.100 ;
        RECT 185.200 86.000 185.600 86.100 ;
        RECT 187.000 86.200 187.400 89.900 ;
        RECT 188.600 87.600 189.000 89.900 ;
        RECT 187.900 87.300 189.000 87.600 ;
        RECT 189.400 87.600 189.800 89.900 ;
        RECT 189.400 87.300 190.500 87.600 ;
        RECT 183.400 85.100 183.700 85.800 ;
        RECT 184.100 85.700 184.500 85.800 ;
        RECT 184.100 85.400 185.800 85.700 ;
        RECT 185.500 85.100 185.800 85.400 ;
        RECT 187.000 85.100 187.300 86.200 ;
        RECT 187.900 85.800 188.200 87.300 ;
        RECT 187.600 85.400 188.200 85.800 ;
        RECT 187.900 85.100 188.200 85.400 ;
        RECT 190.200 85.800 190.500 87.300 ;
        RECT 191.000 86.200 191.400 89.900 ;
        RECT 191.800 87.600 192.200 89.900 ;
        RECT 191.800 87.300 192.900 87.600 ;
        RECT 190.200 85.400 190.800 85.800 ;
        RECT 190.200 85.100 190.500 85.400 ;
        RECT 191.100 85.100 191.400 86.200 ;
        RECT 191.800 85.800 192.200 86.600 ;
        RECT 192.600 85.800 192.900 87.300 ;
        RECT 192.600 85.400 193.200 85.800 ;
        RECT 192.600 85.100 192.900 85.400 ;
        RECT 174.700 84.800 175.200 85.100 ;
        RECT 175.500 84.800 176.200 85.100 ;
        RECT 174.700 82.200 175.100 84.800 ;
        RECT 175.500 84.200 175.800 84.800 ;
        RECT 177.400 84.700 178.300 85.100 ;
        RECT 175.400 83.800 175.800 84.200 ;
        RECT 174.200 81.800 175.100 82.200 ;
        RECT 174.700 81.100 175.100 81.800 ;
        RECT 177.900 82.200 178.300 84.700 ;
        RECT 179.300 84.700 180.200 85.100 ;
        RECT 181.400 84.800 182.600 85.100 ;
        RECT 183.400 84.800 184.400 85.100 ;
        RECT 177.900 81.800 178.600 82.200 ;
        RECT 177.900 81.100 178.300 81.800 ;
        RECT 179.300 81.100 179.700 84.700 ;
        RECT 181.400 81.100 181.800 84.800 ;
        RECT 182.200 84.700 182.600 84.800 ;
        RECT 183.600 81.100 184.400 84.800 ;
        RECT 185.500 84.800 186.600 85.100 ;
        RECT 185.500 84.700 185.900 84.800 ;
        RECT 186.200 81.100 186.600 84.800 ;
        RECT 187.000 81.100 187.400 85.100 ;
        RECT 187.900 84.800 189.000 85.100 ;
        RECT 188.600 81.100 189.000 84.800 ;
        RECT 189.400 84.800 190.500 85.100 ;
        RECT 189.400 81.100 189.800 84.800 ;
        RECT 191.000 81.100 191.400 85.100 ;
        RECT 191.800 84.800 192.900 85.100 ;
        RECT 191.800 81.100 192.200 84.800 ;
        RECT 1.400 75.600 1.800 79.900 ;
        RECT 3.000 75.600 3.400 79.900 ;
        RECT 4.600 75.600 5.000 79.900 ;
        RECT 6.200 75.600 6.600 79.900 ;
        RECT 8.100 76.300 8.500 79.900 ;
        RECT 8.100 75.900 9.000 76.300 ;
        RECT 1.400 75.200 2.300 75.600 ;
        RECT 3.000 75.200 4.100 75.600 ;
        RECT 4.600 75.200 5.700 75.600 ;
        RECT 6.200 75.200 7.400 75.600 ;
        RECT 1.900 74.500 2.300 75.200 ;
        RECT 3.700 74.500 4.100 75.200 ;
        RECT 5.300 74.500 5.700 75.200 ;
        RECT 1.900 74.100 3.200 74.500 ;
        RECT 3.700 74.100 4.900 74.500 ;
        RECT 5.300 74.100 6.600 74.500 ;
        RECT 7.000 74.100 7.400 75.200 ;
        RECT 7.800 74.800 8.200 75.600 ;
        RECT 8.600 75.100 8.900 75.900 ;
        RECT 10.200 75.600 10.600 79.900 ;
        RECT 12.300 77.900 12.900 79.900 ;
        RECT 14.600 77.900 15.000 79.900 ;
        RECT 16.800 78.200 17.200 79.900 ;
        RECT 16.800 77.900 17.800 78.200 ;
        RECT 12.600 77.500 13.000 77.900 ;
        RECT 14.700 77.600 15.000 77.900 ;
        RECT 14.300 77.300 16.100 77.600 ;
        RECT 17.400 77.500 17.800 77.900 ;
        RECT 14.300 77.200 14.700 77.300 ;
        RECT 15.700 77.200 16.100 77.300 ;
        RECT 12.200 76.600 12.900 77.000 ;
        RECT 12.600 76.100 12.900 76.600 ;
        RECT 13.700 76.500 14.800 76.800 ;
        RECT 13.700 76.400 14.100 76.500 ;
        RECT 12.600 75.800 13.800 76.100 ;
        RECT 10.200 75.300 12.300 75.600 ;
        RECT 8.600 74.800 9.700 75.100 ;
        RECT 8.600 74.200 8.900 74.800 ;
        RECT 9.400 74.200 9.700 74.800 ;
        RECT 7.800 74.100 8.200 74.200 ;
        RECT 1.900 73.800 2.300 74.100 ;
        RECT 3.700 73.800 4.100 74.100 ;
        RECT 5.300 73.800 5.700 74.100 ;
        RECT 7.000 73.800 8.200 74.100 ;
        RECT 8.600 73.800 9.000 74.200 ;
        RECT 9.400 73.800 9.800 74.200 ;
        RECT 1.400 73.400 2.300 73.800 ;
        RECT 3.000 73.400 4.100 73.800 ;
        RECT 4.600 73.400 5.700 73.800 ;
        RECT 6.200 73.400 7.400 73.800 ;
        RECT 1.400 71.100 1.800 73.400 ;
        RECT 3.000 71.100 3.400 73.400 ;
        RECT 4.600 71.100 5.000 73.400 ;
        RECT 6.200 71.100 6.600 73.400 ;
        RECT 8.600 72.100 8.900 73.800 ;
        RECT 10.200 73.600 10.600 75.300 ;
        RECT 11.900 75.200 12.300 75.300 ;
        RECT 11.100 74.900 11.500 75.000 ;
        RECT 11.100 74.600 13.000 74.900 ;
        RECT 12.600 74.500 13.000 74.600 ;
        RECT 13.500 74.200 13.800 75.800 ;
        RECT 14.500 75.900 14.800 76.500 ;
        RECT 15.100 76.500 15.500 76.600 ;
        RECT 17.400 76.500 17.800 76.600 ;
        RECT 15.100 76.200 17.800 76.500 ;
        RECT 14.500 75.700 16.900 75.900 ;
        RECT 19.000 75.700 19.400 79.900 ;
        RECT 14.500 75.600 19.400 75.700 ;
        RECT 16.500 75.500 19.400 75.600 ;
        RECT 16.600 75.400 19.400 75.500 ;
        RECT 19.800 75.700 20.200 79.900 ;
        RECT 22.000 78.200 22.400 79.900 ;
        RECT 21.400 77.900 22.400 78.200 ;
        RECT 24.200 77.900 24.600 79.900 ;
        RECT 26.300 77.900 26.900 79.900 ;
        RECT 21.400 77.500 21.800 77.900 ;
        RECT 24.200 77.600 24.500 77.900 ;
        RECT 23.100 77.300 24.900 77.600 ;
        RECT 26.200 77.500 26.600 77.900 ;
        RECT 23.100 77.200 23.500 77.300 ;
        RECT 24.500 77.200 24.900 77.300 ;
        RECT 21.400 76.500 21.800 76.600 ;
        RECT 23.700 76.500 24.100 76.600 ;
        RECT 21.400 76.200 24.100 76.500 ;
        RECT 24.400 76.500 25.500 76.800 ;
        RECT 24.400 75.900 24.700 76.500 ;
        RECT 25.100 76.400 25.500 76.500 ;
        RECT 26.300 76.600 27.000 77.000 ;
        RECT 26.300 76.100 26.600 76.600 ;
        RECT 22.300 75.700 24.700 75.900 ;
        RECT 19.800 75.600 24.700 75.700 ;
        RECT 25.400 75.800 26.600 76.100 ;
        RECT 19.800 75.500 22.700 75.600 ;
        RECT 19.800 75.400 22.600 75.500 ;
        RECT 15.800 75.100 16.200 75.200 ;
        RECT 23.000 75.100 23.400 75.200 ;
        RECT 15.800 74.800 18.300 75.100 ;
        RECT 17.900 74.700 18.300 74.800 ;
        RECT 20.900 74.800 23.400 75.100 ;
        RECT 20.900 74.700 21.300 74.800 ;
        RECT 17.100 74.200 17.500 74.300 ;
        RECT 21.700 74.200 22.100 74.300 ;
        RECT 25.400 74.200 25.700 75.800 ;
        RECT 28.600 75.600 29.000 79.900 ;
        RECT 30.700 76.300 31.100 79.900 ;
        RECT 30.200 75.900 31.100 76.300 ;
        RECT 26.900 75.300 29.000 75.600 ;
        RECT 26.900 75.200 27.300 75.300 ;
        RECT 27.700 74.900 28.100 75.000 ;
        RECT 26.200 74.600 28.100 74.900 ;
        RECT 26.200 74.500 26.600 74.600 ;
        RECT 13.500 74.100 19.000 74.200 ;
        RECT 20.200 74.100 25.700 74.200 ;
        RECT 13.500 73.900 25.700 74.100 ;
        RECT 13.700 73.800 14.100 73.900 ;
        RECT 15.000 73.800 15.400 73.900 ;
        RECT 10.200 73.300 12.100 73.600 ;
        RECT 9.400 72.400 9.800 73.200 ;
        RECT 8.600 71.100 9.000 72.100 ;
        RECT 10.200 71.100 10.600 73.300 ;
        RECT 11.700 73.200 12.100 73.300 ;
        RECT 16.600 72.800 16.900 73.900 ;
        RECT 18.200 73.800 21.000 73.900 ;
        RECT 15.700 72.700 16.100 72.800 ;
        RECT 12.600 72.100 13.000 72.500 ;
        RECT 14.700 72.400 16.100 72.700 ;
        RECT 16.600 72.400 17.000 72.800 ;
        RECT 14.700 72.100 15.000 72.400 ;
        RECT 17.400 72.100 17.800 72.500 ;
        RECT 12.300 71.800 13.000 72.100 ;
        RECT 12.300 71.100 12.900 71.800 ;
        RECT 14.600 71.100 15.000 72.100 ;
        RECT 16.800 71.800 17.800 72.100 ;
        RECT 16.800 71.100 17.200 71.800 ;
        RECT 19.000 71.100 19.400 73.500 ;
        RECT 19.800 71.100 20.200 73.500 ;
        RECT 22.300 72.800 22.600 73.900 ;
        RECT 25.100 73.800 25.500 73.900 ;
        RECT 28.600 73.600 29.000 75.300 ;
        RECT 30.300 74.200 30.600 75.900 ;
        RECT 31.800 75.600 32.200 79.900 ;
        RECT 33.900 77.900 34.500 79.900 ;
        RECT 36.200 77.900 36.600 79.900 ;
        RECT 38.400 78.200 38.800 79.900 ;
        RECT 38.400 77.900 39.400 78.200 ;
        RECT 34.200 77.500 34.600 77.900 ;
        RECT 36.300 77.600 36.600 77.900 ;
        RECT 35.900 77.300 37.700 77.600 ;
        RECT 39.000 77.500 39.400 77.900 ;
        RECT 35.900 77.200 36.300 77.300 ;
        RECT 37.300 77.200 37.700 77.300 ;
        RECT 33.800 76.600 34.500 77.000 ;
        RECT 34.200 76.100 34.500 76.600 ;
        RECT 35.300 76.500 36.400 76.800 ;
        RECT 35.300 76.400 35.700 76.500 ;
        RECT 34.200 75.800 35.400 76.100 ;
        RECT 31.000 74.800 31.400 75.600 ;
        RECT 31.800 75.300 33.900 75.600 ;
        RECT 30.200 73.800 30.600 74.200 ;
        RECT 27.100 73.300 29.000 73.600 ;
        RECT 27.100 73.200 27.500 73.300 ;
        RECT 21.400 72.100 21.800 72.500 ;
        RECT 22.200 72.400 22.600 72.800 ;
        RECT 23.100 72.700 23.500 72.800 ;
        RECT 23.100 72.400 24.500 72.700 ;
        RECT 24.200 72.100 24.500 72.400 ;
        RECT 26.200 72.100 26.600 72.500 ;
        RECT 21.400 71.800 22.400 72.100 ;
        RECT 22.000 71.100 22.400 71.800 ;
        RECT 24.200 71.100 24.600 72.100 ;
        RECT 26.200 71.800 26.900 72.100 ;
        RECT 26.300 71.100 26.900 71.800 ;
        RECT 28.600 71.100 29.000 73.300 ;
        RECT 29.400 72.400 29.800 73.200 ;
        RECT 30.300 72.200 30.600 73.800 ;
        RECT 30.200 71.100 30.600 72.200 ;
        RECT 31.800 73.600 32.200 75.300 ;
        RECT 33.500 75.200 33.900 75.300 ;
        RECT 32.700 74.900 33.100 75.000 ;
        RECT 32.700 74.600 34.600 74.900 ;
        RECT 34.200 74.500 34.600 74.600 ;
        RECT 35.100 74.200 35.400 75.800 ;
        RECT 36.100 75.900 36.400 76.500 ;
        RECT 36.700 76.500 37.100 76.600 ;
        RECT 39.000 76.500 39.400 76.600 ;
        RECT 36.700 76.200 39.400 76.500 ;
        RECT 36.100 75.700 38.500 75.900 ;
        RECT 40.600 75.700 41.000 79.900 ;
        RECT 42.700 79.200 43.100 79.900 ;
        RECT 42.200 78.800 43.100 79.200 ;
        RECT 42.700 76.300 43.100 78.800 ;
        RECT 42.200 75.900 43.100 76.300 ;
        RECT 36.100 75.600 41.000 75.700 ;
        RECT 38.100 75.500 41.000 75.600 ;
        RECT 38.200 75.400 41.000 75.500 ;
        RECT 37.400 75.100 37.800 75.200 ;
        RECT 37.400 74.800 39.900 75.100 ;
        RECT 38.200 74.700 38.600 74.800 ;
        RECT 39.500 74.700 39.900 74.800 ;
        RECT 38.700 74.200 39.100 74.300 ;
        RECT 42.300 74.200 42.600 75.900 ;
        RECT 43.000 74.800 43.400 75.600 ;
        RECT 35.100 73.900 40.600 74.200 ;
        RECT 35.300 73.800 35.700 73.900 ;
        RECT 37.400 73.800 37.800 73.900 ;
        RECT 31.800 73.300 33.700 73.600 ;
        RECT 31.800 71.100 32.200 73.300 ;
        RECT 33.300 73.200 33.700 73.300 ;
        RECT 38.200 72.800 38.500 73.900 ;
        RECT 39.800 73.800 40.600 73.900 ;
        RECT 42.200 73.800 42.600 74.200 ;
        RECT 37.300 72.700 37.700 72.800 ;
        RECT 34.200 72.100 34.600 72.500 ;
        RECT 36.300 72.400 37.700 72.700 ;
        RECT 38.200 72.400 38.600 72.800 ;
        RECT 36.300 72.100 36.600 72.400 ;
        RECT 39.000 72.100 39.400 72.500 ;
        RECT 33.900 71.800 34.600 72.100 ;
        RECT 33.900 71.100 34.500 71.800 ;
        RECT 36.200 71.100 36.600 72.100 ;
        RECT 38.400 71.800 39.400 72.100 ;
        RECT 38.400 71.100 38.800 71.800 ;
        RECT 40.600 71.100 41.000 73.500 ;
        RECT 41.400 72.400 41.800 73.200 ;
        RECT 42.300 72.100 42.600 73.800 ;
        RECT 43.800 73.400 44.200 74.200 ;
        RECT 44.600 73.100 45.000 79.900 ;
        RECT 45.400 75.800 45.800 76.600 ;
        RECT 48.100 76.300 48.500 79.900 ;
        RECT 48.100 75.900 49.000 76.300 ;
        RECT 50.200 76.100 50.600 79.900 ;
        RECT 51.000 76.800 51.400 77.200 ;
        RECT 51.000 76.100 51.300 76.800 ;
        RECT 47.800 74.800 48.200 75.600 ;
        RECT 48.600 75.100 48.900 75.900 ;
        RECT 50.200 75.800 51.300 76.100 ;
        RECT 51.800 75.800 52.200 76.600 ;
        RECT 49.400 75.100 49.800 75.200 ;
        RECT 48.600 74.800 49.800 75.100 ;
        RECT 48.600 74.200 48.900 74.800 ;
        RECT 48.600 73.800 49.000 74.200 ;
        RECT 47.000 73.100 47.400 73.200 ;
        RECT 44.600 72.800 47.400 73.100 ;
        RECT 42.200 71.100 42.600 72.100 ;
        RECT 45.100 71.100 45.500 72.800 ;
        RECT 48.600 72.100 48.900 73.800 ;
        RECT 49.400 72.400 49.800 73.200 ;
        RECT 48.600 71.100 49.000 72.100 ;
        RECT 50.200 71.100 50.600 75.800 ;
        RECT 51.000 72.400 51.400 73.200 ;
        RECT 52.600 73.100 53.000 79.900 ;
        RECT 54.600 76.800 55.000 77.200 ;
        RECT 54.600 76.200 54.900 76.800 ;
        RECT 55.300 76.200 55.700 79.900 ;
        RECT 54.200 75.900 54.900 76.200 ;
        RECT 54.200 75.800 54.600 75.900 ;
        RECT 55.200 75.800 56.200 76.200 ;
        RECT 55.200 74.200 55.500 75.800 ;
        RECT 57.400 75.600 57.800 79.900 ;
        RECT 59.500 79.200 59.900 79.900 ;
        RECT 59.500 78.800 60.200 79.200 ;
        RECT 59.500 76.200 59.900 78.800 ;
        RECT 60.600 76.200 61.000 79.900 ;
        RECT 62.200 76.200 62.600 79.900 ;
        RECT 59.500 75.900 60.200 76.200 ;
        RECT 60.600 75.900 62.600 76.200 ;
        RECT 63.000 75.900 63.400 79.900 ;
        RECT 63.800 77.900 64.200 79.900 ;
        RECT 63.900 77.800 64.200 77.900 ;
        RECT 65.400 77.800 65.800 79.900 ;
        RECT 63.900 77.500 65.700 77.800 ;
        RECT 63.900 76.200 64.200 77.500 ;
        RECT 64.600 76.400 65.000 77.200 ;
        RECT 57.400 75.400 59.400 75.600 ;
        RECT 57.400 75.300 59.500 75.400 ;
        RECT 55.800 74.400 56.200 75.200 ;
        RECT 59.100 75.000 59.500 75.300 ;
        RECT 59.900 75.200 60.200 75.900 ;
        RECT 61.000 75.200 61.400 75.400 ;
        RECT 63.000 75.200 63.300 75.900 ;
        RECT 63.800 75.800 64.200 76.200 ;
        RECT 58.400 74.200 58.800 74.600 ;
        RECT 53.400 73.400 53.800 74.200 ;
        RECT 54.200 73.800 55.500 74.200 ;
        RECT 56.600 74.100 57.000 74.200 ;
        RECT 56.200 73.800 57.700 74.100 ;
        RECT 58.200 73.800 58.700 74.200 ;
        RECT 54.300 73.100 54.600 73.800 ;
        RECT 56.200 73.600 56.600 73.800 ;
        RECT 55.100 73.100 56.900 73.300 ;
        RECT 57.400 73.200 57.700 73.800 ;
        RECT 59.200 73.500 59.500 75.000 ;
        RECT 59.800 74.800 60.200 75.200 ;
        RECT 60.600 74.900 61.400 75.200 ;
        RECT 62.200 74.900 63.400 75.200 ;
        RECT 60.600 74.800 61.000 74.900 ;
        RECT 58.300 73.200 59.500 73.500 ;
        RECT 52.100 72.800 53.000 73.100 ;
        RECT 52.100 72.200 52.500 72.800 ;
        RECT 52.100 71.800 53.000 72.200 ;
        RECT 52.100 71.100 52.500 71.800 ;
        RECT 54.200 71.100 54.600 73.100 ;
        RECT 55.000 73.000 57.000 73.100 ;
        RECT 55.000 71.100 55.400 73.000 ;
        RECT 56.600 71.100 57.000 73.000 ;
        RECT 57.400 72.400 57.800 73.200 ;
        RECT 58.300 72.100 58.600 73.200 ;
        RECT 59.900 73.100 60.200 74.800 ;
        RECT 61.400 73.800 61.800 74.600 ;
        RECT 58.200 71.100 58.600 72.100 ;
        RECT 59.800 71.100 60.200 73.100 ;
        RECT 62.200 73.100 62.500 74.900 ;
        RECT 63.000 74.800 63.400 74.900 ;
        RECT 63.900 74.200 64.200 75.800 ;
        RECT 66.200 75.400 66.600 76.200 ;
        RECT 67.000 75.600 67.400 79.900 ;
        RECT 69.100 77.900 69.700 79.900 ;
        RECT 71.400 77.900 71.800 79.900 ;
        RECT 73.600 78.200 74.000 79.900 ;
        RECT 73.600 77.900 74.600 78.200 ;
        RECT 69.400 77.500 69.800 77.900 ;
        RECT 71.500 77.600 71.800 77.900 ;
        RECT 71.100 77.300 72.900 77.600 ;
        RECT 74.200 77.500 74.600 77.900 ;
        RECT 71.100 77.200 71.500 77.300 ;
        RECT 72.500 77.200 72.900 77.300 ;
        RECT 69.000 76.600 69.700 77.000 ;
        RECT 69.400 76.100 69.700 76.600 ;
        RECT 70.500 76.500 71.600 76.800 ;
        RECT 70.500 76.400 70.900 76.500 ;
        RECT 69.400 75.800 70.600 76.100 ;
        RECT 67.000 75.300 69.100 75.600 ;
        RECT 65.000 74.800 65.800 75.200 ;
        RECT 63.900 74.100 64.700 74.200 ;
        RECT 63.900 73.900 64.800 74.100 ;
        RECT 62.200 71.100 62.600 73.100 ;
        RECT 63.000 72.800 63.400 73.200 ;
        RECT 62.900 72.400 63.300 72.800 ;
        RECT 64.400 71.100 64.800 73.900 ;
        RECT 67.000 73.600 67.400 75.300 ;
        RECT 68.700 75.200 69.100 75.300 ;
        RECT 70.300 75.200 70.600 75.800 ;
        RECT 71.300 75.900 71.600 76.500 ;
        RECT 71.900 76.500 72.300 76.600 ;
        RECT 74.200 76.500 74.600 76.600 ;
        RECT 71.900 76.200 74.600 76.500 ;
        RECT 71.300 75.700 73.700 75.900 ;
        RECT 75.800 75.700 76.200 79.900 ;
        RECT 76.600 76.200 77.000 79.900 ;
        RECT 78.200 76.200 78.600 79.900 ;
        RECT 76.600 75.900 78.600 76.200 ;
        RECT 79.000 75.900 79.400 79.900 ;
        RECT 81.100 76.200 81.500 79.900 ;
        RECT 81.800 76.800 82.200 77.200 ;
        RECT 81.900 76.200 82.200 76.800 ;
        RECT 83.400 76.800 83.800 77.200 ;
        RECT 83.400 76.200 83.700 76.800 ;
        RECT 84.100 76.200 84.500 79.900 ;
        RECT 86.600 76.800 87.000 77.200 ;
        RECT 86.600 76.200 86.900 76.800 ;
        RECT 87.300 76.200 87.700 79.900 ;
        RECT 90.200 76.400 90.600 79.900 ;
        RECT 71.300 75.600 76.200 75.700 ;
        RECT 73.300 75.500 76.200 75.600 ;
        RECT 73.400 75.400 76.200 75.500 ;
        RECT 77.000 75.200 77.400 75.400 ;
        RECT 79.000 75.200 79.300 75.900 ;
        RECT 80.600 75.800 81.600 76.200 ;
        RECT 81.900 76.100 82.600 76.200 ;
        RECT 83.000 76.100 83.700 76.200 ;
        RECT 81.900 75.900 83.700 76.100 ;
        RECT 84.000 75.900 84.500 76.200 ;
        RECT 86.200 75.900 86.900 76.200 ;
        RECT 87.200 75.900 87.700 76.200 ;
        RECT 90.100 75.900 90.600 76.400 ;
        RECT 91.800 76.200 92.200 79.900 ;
        RECT 94.500 76.400 94.900 79.900 ;
        RECT 96.600 77.500 97.000 79.500 ;
        RECT 90.900 75.900 92.200 76.200 ;
        RECT 94.100 76.100 94.900 76.400 ;
        RECT 82.200 75.800 83.400 75.900 ;
        RECT 67.900 74.900 68.300 75.000 ;
        RECT 67.900 74.600 69.800 74.900 ;
        RECT 70.200 74.800 70.600 75.200 ;
        RECT 72.600 75.100 73.000 75.200 ;
        RECT 72.600 74.800 75.100 75.100 ;
        RECT 76.600 74.900 77.400 75.200 ;
        RECT 78.200 74.900 79.400 75.200 ;
        RECT 76.600 74.800 77.000 74.900 ;
        RECT 69.400 74.500 69.800 74.600 ;
        RECT 70.300 74.200 70.600 74.800 ;
        RECT 73.400 74.700 73.800 74.800 ;
        RECT 74.700 74.700 75.100 74.800 ;
        RECT 73.900 74.200 74.300 74.300 ;
        RECT 70.300 73.900 75.800 74.200 ;
        RECT 70.500 73.800 70.900 73.900 ;
        RECT 67.000 73.300 68.900 73.600 ;
        RECT 67.000 71.100 67.400 73.300 ;
        RECT 68.500 73.200 68.900 73.300 ;
        RECT 73.400 72.800 73.700 73.900 ;
        RECT 75.000 73.800 75.800 73.900 ;
        RECT 77.400 73.800 77.800 74.600 ;
        RECT 72.500 72.700 72.900 72.800 ;
        RECT 69.400 72.100 69.800 72.500 ;
        RECT 71.500 72.400 72.900 72.700 ;
        RECT 73.400 72.400 73.800 72.800 ;
        RECT 71.500 72.100 71.800 72.400 ;
        RECT 74.200 72.100 74.600 72.500 ;
        RECT 69.100 71.800 69.800 72.100 ;
        RECT 69.100 71.100 69.700 71.800 ;
        RECT 71.400 71.100 71.800 72.100 ;
        RECT 73.600 71.800 74.600 72.100 ;
        RECT 73.600 71.100 74.000 71.800 ;
        RECT 75.800 71.100 76.200 73.500 ;
        RECT 78.200 73.200 78.500 74.900 ;
        RECT 79.000 74.800 79.400 74.900 ;
        RECT 80.600 74.400 81.000 75.200 ;
        RECT 81.300 74.200 81.600 75.800 ;
        RECT 84.000 74.200 84.300 75.900 ;
        RECT 86.200 75.800 86.600 75.900 ;
        RECT 84.600 74.400 85.000 75.200 ;
        RECT 87.200 74.200 87.500 75.900 ;
        RECT 87.800 74.400 88.200 75.200 ;
        RECT 88.600 74.800 89.000 75.200 ;
        RECT 79.800 74.100 80.200 74.200 ;
        RECT 79.800 73.800 80.600 74.100 ;
        RECT 81.300 73.800 82.600 74.200 ;
        RECT 83.000 73.800 84.300 74.200 ;
        RECT 85.400 74.100 85.800 74.200 ;
        RECT 85.000 73.800 85.800 74.100 ;
        RECT 86.200 73.800 87.500 74.200 ;
        RECT 88.600 74.200 88.900 74.800 ;
        RECT 90.100 74.200 90.400 75.900 ;
        RECT 90.900 74.900 91.200 75.900 ;
        RECT 90.700 74.500 91.200 74.900 ;
        RECT 88.600 74.100 89.000 74.200 ;
        RECT 90.100 74.100 90.600 74.200 ;
        RECT 88.200 73.800 90.600 74.100 ;
        RECT 80.200 73.600 80.600 73.800 ;
        RECT 78.200 71.100 78.600 73.200 ;
        RECT 79.000 72.800 79.400 73.200 ;
        RECT 79.900 73.100 81.700 73.300 ;
        RECT 82.200 73.100 82.500 73.800 ;
        RECT 83.100 73.200 83.400 73.800 ;
        RECT 85.000 73.600 85.400 73.800 ;
        RECT 79.800 73.000 81.800 73.100 ;
        RECT 78.900 72.400 79.300 72.800 ;
        RECT 79.800 71.100 80.200 73.000 ;
        RECT 81.400 71.100 81.800 73.000 ;
        RECT 82.200 71.100 82.600 73.100 ;
        RECT 83.000 71.100 83.400 73.200 ;
        RECT 83.900 73.100 85.700 73.300 ;
        RECT 86.300 73.100 86.600 73.800 ;
        RECT 88.200 73.600 88.600 73.800 ;
        RECT 87.100 73.100 88.900 73.300 ;
        RECT 90.100 73.100 90.400 73.800 ;
        RECT 90.900 73.700 91.200 74.500 ;
        RECT 91.700 74.800 92.200 75.200 ;
        RECT 93.400 74.800 93.800 75.600 ;
        RECT 91.700 74.400 92.100 74.800 ;
        RECT 94.100 74.200 94.400 76.100 ;
        RECT 96.700 75.800 97.000 77.500 ;
        RECT 99.000 76.200 99.400 79.900 ;
        RECT 100.600 76.400 101.000 79.900 ;
        RECT 99.000 75.900 100.300 76.200 ;
        RECT 100.600 75.900 101.100 76.400 ;
        RECT 95.100 75.500 97.000 75.800 ;
        RECT 95.100 74.500 95.400 75.500 ;
        RECT 93.400 73.800 94.400 74.200 ;
        RECT 94.700 74.100 95.400 74.500 ;
        RECT 95.800 74.400 96.200 75.200 ;
        RECT 96.600 74.400 97.000 75.200 ;
        RECT 99.000 74.800 99.500 75.200 ;
        RECT 99.100 74.400 99.500 74.800 ;
        RECT 100.000 74.900 100.300 75.900 ;
        RECT 100.000 74.500 100.500 74.900 ;
        RECT 90.900 73.400 92.200 73.700 ;
        RECT 83.800 73.000 85.800 73.100 ;
        RECT 83.800 71.100 84.200 73.000 ;
        RECT 85.400 71.100 85.800 73.000 ;
        RECT 86.200 71.100 86.600 73.100 ;
        RECT 87.000 73.000 89.000 73.100 ;
        RECT 87.000 71.100 87.400 73.000 ;
        RECT 88.600 71.100 89.000 73.000 ;
        RECT 90.100 72.800 90.600 73.100 ;
        RECT 90.200 71.100 90.600 72.800 ;
        RECT 91.800 71.100 92.200 73.400 ;
        RECT 94.100 73.500 94.400 73.800 ;
        RECT 94.900 73.900 95.400 74.100 ;
        RECT 94.900 73.600 97.000 73.900 ;
        RECT 100.000 73.700 100.300 74.500 ;
        RECT 100.800 74.200 101.100 75.900 ;
        RECT 100.600 73.800 101.100 74.200 ;
        RECT 94.100 73.300 94.500 73.500 ;
        RECT 94.100 73.000 94.900 73.300 ;
        RECT 94.500 72.200 94.900 73.000 ;
        RECT 96.700 72.500 97.000 73.600 ;
        RECT 94.200 71.800 94.900 72.200 ;
        RECT 94.500 71.500 94.900 71.800 ;
        RECT 96.600 71.500 97.000 72.500 ;
        RECT 99.000 73.400 100.300 73.700 ;
        RECT 99.000 71.100 99.400 73.400 ;
        RECT 100.800 73.100 101.100 73.800 ;
        RECT 100.600 72.800 101.100 73.100 ;
        RECT 103.000 75.600 103.400 79.900 ;
        RECT 104.600 75.600 105.000 79.900 ;
        RECT 103.000 75.200 105.000 75.600 ;
        RECT 106.200 75.700 106.600 79.900 ;
        RECT 108.400 78.200 108.800 79.900 ;
        RECT 107.800 77.900 108.800 78.200 ;
        RECT 110.600 77.900 111.000 79.900 ;
        RECT 112.700 77.900 113.300 79.900 ;
        RECT 107.800 77.500 108.200 77.900 ;
        RECT 110.600 77.600 110.900 77.900 ;
        RECT 109.500 77.300 111.300 77.600 ;
        RECT 112.600 77.500 113.000 77.900 ;
        RECT 109.500 77.200 109.900 77.300 ;
        RECT 110.900 77.200 111.300 77.300 ;
        RECT 107.800 76.500 108.200 76.600 ;
        RECT 110.100 76.500 110.500 76.600 ;
        RECT 107.800 76.200 110.500 76.500 ;
        RECT 110.800 76.500 111.900 76.800 ;
        RECT 110.800 75.900 111.100 76.500 ;
        RECT 111.500 76.400 111.900 76.500 ;
        RECT 112.700 76.600 113.400 77.000 ;
        RECT 112.700 76.100 113.000 76.600 ;
        RECT 108.700 75.700 111.100 75.900 ;
        RECT 106.200 75.600 111.100 75.700 ;
        RECT 111.800 75.800 113.000 76.100 ;
        RECT 106.200 75.500 109.100 75.600 ;
        RECT 106.200 75.400 109.000 75.500 ;
        RECT 103.000 73.800 103.400 75.200 ;
        RECT 109.400 75.100 109.800 75.200 ;
        RECT 107.300 74.800 109.800 75.100 ;
        RECT 111.000 75.100 111.400 75.200 ;
        RECT 111.800 75.100 112.100 75.800 ;
        RECT 115.000 75.600 115.400 79.900 ;
        RECT 113.300 75.300 115.400 75.600 ;
        RECT 115.800 75.700 116.200 79.900 ;
        RECT 118.000 78.200 118.400 79.900 ;
        RECT 117.400 77.900 118.400 78.200 ;
        RECT 120.200 77.900 120.600 79.900 ;
        RECT 122.300 77.900 122.900 79.900 ;
        RECT 117.400 77.500 117.800 77.900 ;
        RECT 120.200 77.600 120.500 77.900 ;
        RECT 119.100 77.300 120.900 77.600 ;
        RECT 122.200 77.500 122.600 77.900 ;
        RECT 119.100 77.200 119.500 77.300 ;
        RECT 120.500 77.200 120.900 77.300 ;
        RECT 117.400 76.500 117.800 76.600 ;
        RECT 119.700 76.500 120.100 76.600 ;
        RECT 117.400 76.200 120.100 76.500 ;
        RECT 120.400 76.500 121.500 76.800 ;
        RECT 120.400 75.900 120.700 76.500 ;
        RECT 121.100 76.400 121.500 76.500 ;
        RECT 122.300 76.600 123.000 77.000 ;
        RECT 122.300 76.100 122.600 76.600 ;
        RECT 118.300 75.700 120.700 75.900 ;
        RECT 115.800 75.600 120.700 75.700 ;
        RECT 121.400 75.800 122.600 76.100 ;
        RECT 115.800 75.500 118.700 75.600 ;
        RECT 115.800 75.400 118.600 75.500 ;
        RECT 113.300 75.200 113.700 75.300 ;
        RECT 111.000 74.800 112.100 75.100 ;
        RECT 114.100 74.900 114.500 75.000 ;
        RECT 107.300 74.700 107.700 74.800 ;
        RECT 108.100 74.200 108.500 74.300 ;
        RECT 111.800 74.200 112.100 74.800 ;
        RECT 112.600 74.600 114.500 74.900 ;
        RECT 112.600 74.500 113.000 74.600 ;
        RECT 103.000 73.400 105.000 73.800 ;
        RECT 105.400 73.400 105.800 74.200 ;
        RECT 106.600 73.900 112.100 74.200 ;
        RECT 106.600 73.800 107.400 73.900 ;
        RECT 100.600 71.100 101.000 72.800 ;
        RECT 103.000 71.100 103.400 73.400 ;
        RECT 104.600 71.100 105.000 73.400 ;
        RECT 106.200 71.100 106.600 73.500 ;
        RECT 108.700 72.800 109.000 73.900 ;
        RECT 111.500 73.800 111.900 73.900 ;
        RECT 115.000 73.600 115.400 75.300 ;
        RECT 121.400 75.200 121.700 75.800 ;
        RECT 123.000 75.600 123.400 76.200 ;
        RECT 124.600 75.600 125.000 79.900 ;
        RECT 125.700 76.300 126.100 79.900 ;
        RECT 125.700 75.900 126.600 76.300 ;
        RECT 122.900 75.300 125.000 75.600 ;
        RECT 122.900 75.200 123.300 75.300 ;
        RECT 119.000 75.100 119.400 75.200 ;
        RECT 116.900 74.800 119.400 75.100 ;
        RECT 121.400 74.800 121.800 75.200 ;
        RECT 123.700 74.900 124.100 75.000 ;
        RECT 116.900 74.700 117.300 74.800 ;
        RECT 117.700 74.200 118.100 74.300 ;
        RECT 121.400 74.200 121.700 74.800 ;
        RECT 122.200 74.600 124.100 74.900 ;
        RECT 122.200 74.500 122.600 74.600 ;
        RECT 116.200 73.900 121.700 74.200 ;
        RECT 116.200 73.800 117.000 73.900 ;
        RECT 113.500 73.300 115.400 73.600 ;
        RECT 113.500 73.200 113.900 73.300 ;
        RECT 107.800 72.100 108.200 72.500 ;
        RECT 108.600 72.400 109.000 72.800 ;
        RECT 109.500 72.700 109.900 72.800 ;
        RECT 109.500 72.400 110.900 72.700 ;
        RECT 110.600 72.100 110.900 72.400 ;
        RECT 112.600 72.100 113.000 72.500 ;
        RECT 107.800 71.800 108.800 72.100 ;
        RECT 108.400 71.100 108.800 71.800 ;
        RECT 110.600 71.100 111.000 72.100 ;
        RECT 112.600 71.800 113.300 72.100 ;
        RECT 112.700 71.100 113.300 71.800 ;
        RECT 115.000 71.100 115.400 73.300 ;
        RECT 115.800 71.100 116.200 73.500 ;
        RECT 118.300 72.800 118.600 73.900 ;
        RECT 121.100 73.800 121.500 73.900 ;
        RECT 124.600 73.600 125.000 75.300 ;
        RECT 125.400 74.800 125.800 75.600 ;
        RECT 126.200 74.200 126.500 75.900 ;
        RECT 128.600 75.600 129.000 79.900 ;
        RECT 130.200 75.600 130.600 79.900 ;
        RECT 131.800 75.600 132.200 79.900 ;
        RECT 133.400 75.600 133.800 79.900 ;
        RECT 135.800 75.600 136.200 79.900 ;
        RECT 137.400 75.600 137.800 79.900 ;
        RECT 128.600 75.200 129.500 75.600 ;
        RECT 130.200 75.200 131.300 75.600 ;
        RECT 131.800 75.200 132.900 75.600 ;
        RECT 133.400 75.200 134.600 75.600 ;
        RECT 129.100 74.500 129.500 75.200 ;
        RECT 130.900 74.500 131.300 75.200 ;
        RECT 132.500 74.500 132.900 75.200 ;
        RECT 123.100 73.300 125.000 73.600 ;
        RECT 123.100 73.200 123.500 73.300 ;
        RECT 117.400 72.100 117.800 72.500 ;
        RECT 118.200 72.400 118.600 72.800 ;
        RECT 119.100 72.700 119.500 72.800 ;
        RECT 119.100 72.400 120.500 72.700 ;
        RECT 120.200 72.100 120.500 72.400 ;
        RECT 122.200 72.100 122.600 72.500 ;
        RECT 117.400 71.800 118.400 72.100 ;
        RECT 118.000 71.100 118.400 71.800 ;
        RECT 120.200 71.100 120.600 72.100 ;
        RECT 122.200 71.800 122.900 72.100 ;
        RECT 122.300 71.100 122.900 71.800 ;
        RECT 124.600 71.100 125.000 73.300 ;
        RECT 125.400 73.800 125.800 74.200 ;
        RECT 126.200 73.800 126.600 74.200 ;
        RECT 129.100 74.100 130.400 74.500 ;
        RECT 130.900 74.100 132.100 74.500 ;
        RECT 132.500 74.100 133.800 74.500 ;
        RECT 134.200 74.100 134.600 75.200 ;
        RECT 135.800 75.200 137.800 75.600 ;
        RECT 139.000 75.700 139.400 79.900 ;
        RECT 141.200 78.200 141.600 79.900 ;
        RECT 140.600 77.900 141.600 78.200 ;
        RECT 143.400 77.900 143.800 79.900 ;
        RECT 145.500 77.900 146.100 79.900 ;
        RECT 140.600 77.500 141.000 77.900 ;
        RECT 143.400 77.600 143.700 77.900 ;
        RECT 142.300 77.300 144.100 77.600 ;
        RECT 145.400 77.500 145.800 77.900 ;
        RECT 142.300 77.200 142.700 77.300 ;
        RECT 143.700 77.200 144.100 77.300 ;
        RECT 140.600 76.500 141.000 76.600 ;
        RECT 142.900 76.500 143.300 76.600 ;
        RECT 140.600 76.200 143.300 76.500 ;
        RECT 143.600 76.500 144.700 76.800 ;
        RECT 143.600 75.900 143.900 76.500 ;
        RECT 144.300 76.400 144.700 76.500 ;
        RECT 145.500 76.600 146.200 77.000 ;
        RECT 145.500 76.100 145.800 76.600 ;
        RECT 141.500 75.700 143.900 75.900 ;
        RECT 139.000 75.600 143.900 75.700 ;
        RECT 144.600 75.800 145.800 76.100 ;
        RECT 139.000 75.500 141.900 75.600 ;
        RECT 139.000 75.400 141.800 75.500 ;
        RECT 135.000 74.100 135.400 74.200 ;
        RECT 129.100 73.800 129.500 74.100 ;
        RECT 130.900 73.800 131.300 74.100 ;
        RECT 132.500 73.800 132.900 74.100 ;
        RECT 134.200 73.800 135.400 74.100 ;
        RECT 135.800 73.800 136.200 75.200 ;
        RECT 142.200 75.100 142.600 75.200 ;
        RECT 140.100 74.800 142.600 75.100 ;
        RECT 140.100 74.700 140.500 74.800 ;
        RECT 140.900 74.200 141.300 74.300 ;
        RECT 144.600 74.200 144.900 75.800 ;
        RECT 147.800 75.600 148.200 79.900 ;
        RECT 150.200 76.200 150.600 79.900 ;
        RECT 150.200 75.900 151.300 76.200 ;
        RECT 151.800 75.900 152.200 79.900 ;
        RECT 146.100 75.300 148.200 75.600 ;
        RECT 146.100 75.200 146.500 75.300 ;
        RECT 146.900 74.900 147.300 75.000 ;
        RECT 145.400 74.600 147.300 74.900 ;
        RECT 145.400 74.500 145.800 74.600 ;
        RECT 138.200 74.100 138.600 74.200 ;
        RECT 139.400 74.100 144.900 74.200 ;
        RECT 138.200 73.900 144.900 74.100 ;
        RECT 138.200 73.800 140.200 73.900 ;
        RECT 125.400 73.100 125.700 73.800 ;
        RECT 126.200 73.100 126.500 73.800 ;
        RECT 128.600 73.400 129.500 73.800 ;
        RECT 130.200 73.400 131.300 73.800 ;
        RECT 131.800 73.400 132.900 73.800 ;
        RECT 133.400 73.400 134.600 73.800 ;
        RECT 135.800 73.400 137.800 73.800 ;
        RECT 138.200 73.400 138.600 73.800 ;
        RECT 125.400 72.800 126.500 73.100 ;
        RECT 126.200 72.100 126.500 72.800 ;
        RECT 127.000 72.400 127.400 73.200 ;
        RECT 126.200 71.100 126.600 72.100 ;
        RECT 128.600 71.100 129.000 73.400 ;
        RECT 130.200 71.100 130.600 73.400 ;
        RECT 131.800 71.100 132.200 73.400 ;
        RECT 133.400 71.100 133.800 73.400 ;
        RECT 135.800 71.100 136.200 73.400 ;
        RECT 137.400 71.100 137.800 73.400 ;
        RECT 139.000 71.100 139.400 73.500 ;
        RECT 141.500 72.800 141.800 73.900 ;
        RECT 144.300 73.800 144.700 73.900 ;
        RECT 147.800 73.600 148.200 75.300 ;
        RECT 151.000 75.600 151.300 75.900 ;
        RECT 151.000 75.200 151.600 75.600 ;
        RECT 151.000 73.700 151.300 75.200 ;
        RECT 151.900 74.800 152.200 75.900 ;
        RECT 146.300 73.300 148.200 73.600 ;
        RECT 146.300 73.200 146.700 73.300 ;
        RECT 140.600 72.100 141.000 72.500 ;
        RECT 141.400 72.400 141.800 72.800 ;
        RECT 142.300 72.700 142.700 72.800 ;
        RECT 142.300 72.400 143.700 72.700 ;
        RECT 143.400 72.100 143.700 72.400 ;
        RECT 145.400 72.100 145.800 72.500 ;
        RECT 140.600 71.800 141.600 72.100 ;
        RECT 141.200 71.100 141.600 71.800 ;
        RECT 143.400 71.100 143.800 72.100 ;
        RECT 145.400 71.800 146.100 72.100 ;
        RECT 145.500 71.100 146.100 71.800 ;
        RECT 147.800 71.100 148.200 73.300 ;
        RECT 150.200 73.400 151.300 73.700 ;
        RECT 150.200 71.100 150.600 73.400 ;
        RECT 151.800 71.100 152.200 74.800 ;
        RECT 152.600 72.400 153.000 73.200 ;
        RECT 153.400 71.100 153.800 79.900 ;
        RECT 154.200 75.700 154.600 79.900 ;
        RECT 156.400 78.200 156.800 79.900 ;
        RECT 155.800 77.900 156.800 78.200 ;
        RECT 158.600 77.900 159.000 79.900 ;
        RECT 160.700 77.900 161.300 79.900 ;
        RECT 155.800 77.500 156.200 77.900 ;
        RECT 158.600 77.600 158.900 77.900 ;
        RECT 157.500 77.300 159.300 77.600 ;
        RECT 160.600 77.500 161.000 77.900 ;
        RECT 157.500 77.200 157.900 77.300 ;
        RECT 158.900 77.200 159.300 77.300 ;
        RECT 155.800 76.500 156.200 76.600 ;
        RECT 158.100 76.500 158.500 76.600 ;
        RECT 155.800 76.200 158.500 76.500 ;
        RECT 158.800 76.500 159.900 76.800 ;
        RECT 158.800 75.900 159.100 76.500 ;
        RECT 159.500 76.400 159.900 76.500 ;
        RECT 160.700 76.600 161.400 77.000 ;
        RECT 160.700 76.100 161.000 76.600 ;
        RECT 156.700 75.700 159.100 75.900 ;
        RECT 154.200 75.600 159.100 75.700 ;
        RECT 159.800 75.800 161.000 76.100 ;
        RECT 154.200 75.500 157.100 75.600 ;
        RECT 154.200 75.400 157.000 75.500 ;
        RECT 157.400 75.100 157.800 75.200 ;
        RECT 158.200 75.100 158.600 75.200 ;
        RECT 155.300 74.800 158.600 75.100 ;
        RECT 155.300 74.700 155.700 74.800 ;
        RECT 156.100 74.200 156.500 74.300 ;
        RECT 159.800 74.200 160.100 75.800 ;
        RECT 163.000 75.600 163.400 79.900 ;
        RECT 164.100 76.300 164.500 79.900 ;
        RECT 164.100 75.900 165.000 76.300 ;
        RECT 161.300 75.300 163.400 75.600 ;
        RECT 161.300 75.200 161.700 75.300 ;
        RECT 162.100 74.900 162.500 75.000 ;
        RECT 160.600 74.600 162.500 74.900 ;
        RECT 160.600 74.500 161.000 74.600 ;
        RECT 154.600 73.900 160.100 74.200 ;
        RECT 154.600 73.800 155.400 73.900 ;
        RECT 154.200 71.100 154.600 73.500 ;
        RECT 156.700 72.800 157.000 73.900 ;
        RECT 159.500 73.800 159.900 73.900 ;
        RECT 163.000 73.600 163.400 75.300 ;
        RECT 163.800 74.800 164.200 75.600 ;
        RECT 164.600 75.100 164.900 75.900 ;
        RECT 165.400 75.100 165.800 75.200 ;
        RECT 164.600 74.800 165.800 75.100 ;
        RECT 161.500 73.300 163.400 73.600 ;
        RECT 161.500 73.200 161.900 73.300 ;
        RECT 155.800 72.100 156.200 72.500 ;
        RECT 156.600 72.400 157.000 72.800 ;
        RECT 157.500 72.700 157.900 72.800 ;
        RECT 157.500 72.400 158.900 72.700 ;
        RECT 158.600 72.100 158.900 72.400 ;
        RECT 160.600 72.100 161.000 72.500 ;
        RECT 155.800 71.800 156.800 72.100 ;
        RECT 156.400 71.100 156.800 71.800 ;
        RECT 158.600 71.100 159.000 72.100 ;
        RECT 160.600 71.800 161.300 72.100 ;
        RECT 160.700 71.100 161.300 71.800 ;
        RECT 163.000 71.100 163.400 73.300 ;
        RECT 164.600 74.200 164.900 74.800 ;
        RECT 164.600 73.800 165.000 74.200 ;
        RECT 164.600 72.100 164.900 73.800 ;
        RECT 166.200 73.400 166.600 74.200 ;
        RECT 165.400 72.400 165.800 73.200 ;
        RECT 167.000 73.100 167.400 79.900 ;
        RECT 167.800 75.800 168.200 76.600 ;
        RECT 169.400 76.100 169.800 79.900 ;
        RECT 170.600 76.800 171.000 77.200 ;
        RECT 170.600 76.200 170.900 76.800 ;
        RECT 171.300 76.200 171.700 79.900 ;
        RECT 170.200 76.100 170.900 76.200 ;
        RECT 169.400 75.900 170.900 76.100 ;
        RECT 171.200 75.900 171.700 76.200 ;
        RECT 169.400 75.800 170.600 75.900 ;
        RECT 167.000 72.800 167.900 73.100 ;
        RECT 167.500 72.200 167.900 72.800 ;
        RECT 168.600 72.400 169.000 73.200 ;
        RECT 164.600 71.100 165.000 72.100 ;
        RECT 167.000 71.800 167.900 72.200 ;
        RECT 167.500 71.100 167.900 71.800 ;
        RECT 169.400 71.100 169.800 75.800 ;
        RECT 170.200 75.100 170.600 75.200 ;
        RECT 171.200 75.100 171.500 75.900 ;
        RECT 170.200 74.800 171.500 75.100 ;
        RECT 171.200 74.200 171.500 74.800 ;
        RECT 171.800 75.100 172.200 75.200 ;
        RECT 174.200 75.100 174.600 79.900 ;
        RECT 175.300 76.300 175.700 79.900 ;
        RECT 175.300 75.900 176.200 76.300 ;
        RECT 177.400 75.900 177.800 79.900 ;
        RECT 178.200 76.200 178.600 79.900 ;
        RECT 179.800 76.200 180.200 79.900 ;
        RECT 178.200 75.900 180.200 76.200 ;
        RECT 175.000 75.100 175.400 75.600 ;
        RECT 171.800 74.800 175.400 75.100 ;
        RECT 171.800 74.400 172.200 74.800 ;
        RECT 170.200 73.800 171.500 74.200 ;
        RECT 172.600 74.100 173.000 74.200 ;
        RECT 172.200 73.800 173.000 74.100 ;
        RECT 170.300 73.100 170.600 73.800 ;
        RECT 172.200 73.600 172.600 73.800 ;
        RECT 171.100 73.100 172.900 73.300 ;
        RECT 170.200 71.100 170.600 73.100 ;
        RECT 171.000 73.000 173.000 73.100 ;
        RECT 171.000 71.100 171.400 73.000 ;
        RECT 172.600 71.100 173.000 73.000 ;
        RECT 173.400 72.400 173.800 73.200 ;
        RECT 174.200 71.100 174.600 74.800 ;
        RECT 175.800 74.200 176.100 75.900 ;
        RECT 177.500 75.200 177.800 75.900 ;
        RECT 180.600 75.800 181.000 76.600 ;
        RECT 179.400 75.200 179.800 75.400 ;
        RECT 177.400 74.900 178.600 75.200 ;
        RECT 179.400 74.900 180.200 75.200 ;
        RECT 177.400 74.800 177.800 74.900 ;
        RECT 175.800 73.800 176.200 74.200 ;
        RECT 175.800 72.200 176.100 73.800 ;
        RECT 176.600 72.400 177.000 73.200 ;
        RECT 177.400 72.800 177.800 73.200 ;
        RECT 178.300 73.100 178.600 74.900 ;
        RECT 179.800 74.800 180.200 74.900 ;
        RECT 179.000 74.100 179.400 74.600 ;
        RECT 181.400 74.100 181.800 79.900 ;
        RECT 179.000 73.800 181.800 74.100 ;
        RECT 181.400 73.100 181.800 73.800 ;
        RECT 182.200 74.100 182.600 74.200 ;
        RECT 183.000 74.100 183.400 79.900 ;
        RECT 184.600 75.700 185.000 79.900 ;
        RECT 186.800 78.200 187.200 79.900 ;
        RECT 186.200 77.900 187.200 78.200 ;
        RECT 189.000 77.900 189.400 79.900 ;
        RECT 191.100 77.900 191.700 79.900 ;
        RECT 186.200 77.500 186.600 77.900 ;
        RECT 189.000 77.600 189.300 77.900 ;
        RECT 187.900 77.300 189.700 77.600 ;
        RECT 191.000 77.500 191.400 77.900 ;
        RECT 187.900 77.200 188.300 77.300 ;
        RECT 189.300 77.200 189.700 77.300 ;
        RECT 186.200 76.500 186.600 76.600 ;
        RECT 188.500 76.500 188.900 76.600 ;
        RECT 186.200 76.200 188.900 76.500 ;
        RECT 189.200 76.500 190.300 76.800 ;
        RECT 189.200 75.900 189.500 76.500 ;
        RECT 189.900 76.400 190.300 76.500 ;
        RECT 191.100 76.600 191.800 77.000 ;
        RECT 191.100 76.100 191.400 76.600 ;
        RECT 187.100 75.700 189.500 75.900 ;
        RECT 184.600 75.600 189.500 75.700 ;
        RECT 190.200 75.800 191.400 76.100 ;
        RECT 184.600 75.500 187.500 75.600 ;
        RECT 184.600 75.400 187.400 75.500 ;
        RECT 187.800 75.100 188.200 75.200 ;
        RECT 185.700 74.800 188.200 75.100 ;
        RECT 185.700 74.700 186.100 74.800 ;
        RECT 187.000 74.700 187.400 74.800 ;
        RECT 186.500 74.200 186.900 74.300 ;
        RECT 190.200 74.200 190.500 75.800 ;
        RECT 193.400 75.600 193.800 79.900 ;
        RECT 191.700 75.300 193.800 75.600 ;
        RECT 191.700 75.200 192.100 75.300 ;
        RECT 192.500 74.900 192.900 75.000 ;
        RECT 191.000 74.600 192.900 74.900 ;
        RECT 191.000 74.500 191.400 74.600 ;
        RECT 182.200 73.800 183.400 74.100 ;
        RECT 185.000 73.900 190.500 74.200 ;
        RECT 185.000 73.800 185.800 73.900 ;
        RECT 182.200 73.400 182.600 73.800 ;
        RECT 177.500 72.400 177.900 72.800 ;
        RECT 175.800 71.100 176.200 72.200 ;
        RECT 178.200 71.100 178.600 73.100 ;
        RECT 180.900 72.800 181.800 73.100 ;
        RECT 180.900 71.100 181.300 72.800 ;
        RECT 183.000 71.100 183.400 73.800 ;
        RECT 183.800 72.400 184.200 73.200 ;
        RECT 184.600 71.100 185.000 73.500 ;
        RECT 187.100 72.800 187.400 73.900 ;
        RECT 189.900 73.800 190.300 73.900 ;
        RECT 193.400 73.600 193.800 75.300 ;
        RECT 191.900 73.300 193.800 73.600 ;
        RECT 191.900 73.200 192.300 73.300 ;
        RECT 186.200 72.100 186.600 72.500 ;
        RECT 187.000 72.400 187.400 72.800 ;
        RECT 187.900 72.700 188.300 72.800 ;
        RECT 187.900 72.400 189.300 72.700 ;
        RECT 189.000 72.100 189.300 72.400 ;
        RECT 191.000 72.100 191.400 72.500 ;
        RECT 186.200 71.800 187.200 72.100 ;
        RECT 186.800 71.100 187.200 71.800 ;
        RECT 189.000 71.100 189.400 72.100 ;
        RECT 191.000 71.800 191.700 72.100 ;
        RECT 191.100 71.100 191.700 71.800 ;
        RECT 193.400 71.100 193.800 73.300 ;
        RECT 2.200 67.600 2.600 69.900 ;
        RECT 1.500 67.300 2.600 67.600 ;
        RECT 3.800 67.600 4.200 69.900 ;
        RECT 5.400 67.600 5.800 69.900 ;
        RECT 7.000 67.600 7.400 69.900 ;
        RECT 8.600 67.600 9.000 69.900 ;
        RECT 10.200 67.700 10.600 69.900 ;
        RECT 12.300 69.200 12.900 69.900 ;
        RECT 12.300 68.900 13.000 69.200 ;
        RECT 14.600 68.900 15.000 69.900 ;
        RECT 16.800 69.200 17.200 69.900 ;
        RECT 16.800 68.900 17.800 69.200 ;
        RECT 12.600 68.500 13.000 68.900 ;
        RECT 14.700 68.600 15.000 68.900 ;
        RECT 14.700 68.300 16.100 68.600 ;
        RECT 15.700 68.200 16.100 68.300 ;
        RECT 16.600 68.200 17.000 68.600 ;
        RECT 17.400 68.500 17.800 68.900 ;
        RECT 11.700 67.700 12.100 67.800 ;
        RECT 1.500 65.800 1.800 67.300 ;
        RECT 3.800 67.200 4.700 67.600 ;
        RECT 5.400 67.200 6.500 67.600 ;
        RECT 7.000 67.200 8.100 67.600 ;
        RECT 8.600 67.200 9.800 67.600 ;
        RECT 4.300 66.900 4.700 67.200 ;
        RECT 6.100 66.900 6.500 67.200 ;
        RECT 7.700 66.900 8.100 67.200 ;
        RECT 4.300 66.500 5.600 66.900 ;
        RECT 6.100 66.500 7.300 66.900 ;
        RECT 7.700 66.500 9.000 66.900 ;
        RECT 4.300 65.800 4.700 66.500 ;
        RECT 6.100 65.800 6.500 66.500 ;
        RECT 7.700 65.800 8.100 66.500 ;
        RECT 9.400 65.800 9.800 67.200 ;
        RECT 1.200 65.400 1.800 65.800 ;
        RECT 1.500 65.100 1.800 65.400 ;
        RECT 3.800 65.400 4.700 65.800 ;
        RECT 5.400 65.400 6.500 65.800 ;
        RECT 7.000 65.400 8.100 65.800 ;
        RECT 8.600 65.400 9.800 65.800 ;
        RECT 10.200 67.400 12.100 67.700 ;
        RECT 10.200 65.700 10.600 67.400 ;
        RECT 13.700 67.100 14.100 67.200 ;
        RECT 16.600 67.100 16.900 68.200 ;
        RECT 19.000 67.500 19.400 69.900 ;
        RECT 19.800 67.900 20.200 69.900 ;
        RECT 20.600 68.000 21.000 69.900 ;
        RECT 22.200 68.000 22.600 69.900 ;
        RECT 20.600 67.900 22.600 68.000 ;
        RECT 19.900 67.200 20.200 67.900 ;
        RECT 20.700 67.700 22.500 67.900 ;
        RECT 21.800 67.200 22.200 67.400 ;
        RECT 18.200 67.100 19.000 67.200 ;
        RECT 13.500 66.800 19.000 67.100 ;
        RECT 19.800 66.800 21.100 67.200 ;
        RECT 21.800 67.100 22.600 67.200 ;
        RECT 23.000 67.100 23.400 69.900 ;
        RECT 23.800 67.800 24.200 68.600 ;
        RECT 24.600 67.500 25.000 69.900 ;
        RECT 26.800 69.200 27.200 69.900 ;
        RECT 26.200 68.900 27.200 69.200 ;
        RECT 29.000 68.900 29.400 69.900 ;
        RECT 31.100 69.200 31.700 69.900 ;
        RECT 31.000 68.900 31.700 69.200 ;
        RECT 26.200 68.500 26.600 68.900 ;
        RECT 29.000 68.600 29.300 68.900 ;
        RECT 27.000 68.200 27.400 68.600 ;
        RECT 27.900 68.300 29.300 68.600 ;
        RECT 31.000 68.500 31.400 68.900 ;
        RECT 27.900 68.200 28.300 68.300 ;
        RECT 27.100 67.200 27.400 68.200 ;
        RECT 31.900 67.700 32.300 67.800 ;
        RECT 33.400 67.700 33.800 69.900 ;
        RECT 34.200 67.900 34.600 69.900 ;
        RECT 35.000 68.000 35.400 69.900 ;
        RECT 36.600 68.000 37.000 69.900 ;
        RECT 35.000 67.900 37.000 68.000 ;
        RECT 31.900 67.400 33.800 67.700 ;
        RECT 21.800 66.900 23.400 67.100 ;
        RECT 22.200 66.800 23.400 66.900 ;
        RECT 25.000 67.100 25.800 67.200 ;
        RECT 27.000 67.100 27.400 67.200 ;
        RECT 29.900 67.100 30.300 67.200 ;
        RECT 25.000 66.800 30.500 67.100 ;
        RECT 12.600 66.400 13.000 66.500 ;
        RECT 11.100 66.100 13.000 66.400 ;
        RECT 11.100 66.000 11.500 66.100 ;
        RECT 11.900 65.700 12.300 65.800 ;
        RECT 10.200 65.400 12.300 65.700 ;
        RECT 1.500 64.800 2.600 65.100 ;
        RECT 2.200 61.100 2.600 64.800 ;
        RECT 3.800 61.100 4.200 65.400 ;
        RECT 5.400 61.100 5.800 65.400 ;
        RECT 7.000 61.100 7.400 65.400 ;
        RECT 8.600 61.100 9.000 65.400 ;
        RECT 10.200 61.100 10.600 65.400 ;
        RECT 13.500 65.200 13.800 66.800 ;
        RECT 17.100 66.700 17.500 66.800 ;
        RECT 16.600 66.200 17.000 66.300 ;
        RECT 17.900 66.200 18.300 66.300 ;
        RECT 15.800 65.900 18.300 66.200 ;
        RECT 15.800 65.800 16.200 65.900 ;
        RECT 16.600 65.500 19.400 65.600 ;
        RECT 16.500 65.400 19.400 65.500 ;
        RECT 12.600 64.900 13.800 65.200 ;
        RECT 14.500 65.300 19.400 65.400 ;
        RECT 14.500 65.100 16.900 65.300 ;
        RECT 12.600 64.400 12.900 64.900 ;
        RECT 12.200 64.000 12.900 64.400 ;
        RECT 13.700 64.500 14.100 64.600 ;
        RECT 14.500 64.500 14.800 65.100 ;
        RECT 13.700 64.200 14.800 64.500 ;
        RECT 15.100 64.500 17.800 64.800 ;
        RECT 15.100 64.400 15.500 64.500 ;
        RECT 17.400 64.400 17.800 64.500 ;
        RECT 14.300 63.700 14.700 63.800 ;
        RECT 15.700 63.700 16.100 63.800 ;
        RECT 12.600 63.100 13.000 63.500 ;
        RECT 14.300 63.400 16.100 63.700 ;
        RECT 14.700 63.100 15.000 63.400 ;
        RECT 17.400 63.100 17.800 63.500 ;
        RECT 12.300 61.100 12.900 63.100 ;
        RECT 14.600 61.100 15.000 63.100 ;
        RECT 16.800 62.800 17.800 63.100 ;
        RECT 16.800 61.100 17.200 62.800 ;
        RECT 19.000 61.100 19.400 65.300 ;
        RECT 19.800 65.100 20.200 65.200 ;
        RECT 20.800 65.100 21.100 66.800 ;
        RECT 21.400 66.100 21.800 66.600 ;
        RECT 22.200 66.100 22.600 66.200 ;
        RECT 21.400 65.800 22.600 66.100 ;
        RECT 19.800 64.800 20.500 65.100 ;
        RECT 20.800 64.800 21.300 65.100 ;
        RECT 20.200 64.200 20.500 64.800 ;
        RECT 20.200 63.800 20.600 64.200 ;
        RECT 20.900 61.100 21.300 64.800 ;
        RECT 23.000 61.100 23.400 66.800 ;
        RECT 26.500 66.700 26.900 66.800 ;
        RECT 25.700 66.200 26.100 66.300 ;
        RECT 25.700 66.100 28.200 66.200 ;
        RECT 29.400 66.100 29.800 66.200 ;
        RECT 25.700 65.900 29.800 66.100 ;
        RECT 27.800 65.800 29.800 65.900 ;
        RECT 24.600 65.500 27.400 65.600 ;
        RECT 24.600 65.400 27.500 65.500 ;
        RECT 24.600 65.300 29.500 65.400 ;
        RECT 24.600 61.100 25.000 65.300 ;
        RECT 27.100 65.100 29.500 65.300 ;
        RECT 26.200 64.500 28.900 64.800 ;
        RECT 26.200 64.400 26.600 64.500 ;
        RECT 28.500 64.400 28.900 64.500 ;
        RECT 29.200 64.500 29.500 65.100 ;
        RECT 30.200 65.200 30.500 66.800 ;
        RECT 31.000 66.400 31.400 66.500 ;
        RECT 31.000 66.100 32.900 66.400 ;
        RECT 32.500 66.000 32.900 66.100 ;
        RECT 31.700 65.700 32.100 65.800 ;
        RECT 33.400 65.700 33.800 67.400 ;
        RECT 34.300 67.200 34.600 67.900 ;
        RECT 35.100 67.700 36.900 67.900 ;
        RECT 36.200 67.200 36.600 67.400 ;
        RECT 34.200 66.800 35.500 67.200 ;
        RECT 36.200 67.100 37.000 67.200 ;
        RECT 37.400 67.100 37.800 69.900 ;
        RECT 38.200 67.800 38.600 68.600 ;
        RECT 39.000 67.500 39.400 69.900 ;
        RECT 41.200 69.200 41.600 69.900 ;
        RECT 40.600 68.900 41.600 69.200 ;
        RECT 43.400 68.900 43.800 69.900 ;
        RECT 45.500 69.200 46.100 69.900 ;
        RECT 45.400 68.900 46.100 69.200 ;
        RECT 47.800 69.100 48.200 69.900 ;
        RECT 48.600 69.100 49.000 69.200 ;
        RECT 40.600 68.500 41.000 68.900 ;
        RECT 43.400 68.600 43.700 68.900 ;
        RECT 41.400 68.200 41.800 68.600 ;
        RECT 42.300 68.300 43.700 68.600 ;
        RECT 45.400 68.500 45.800 68.900 ;
        RECT 47.800 68.800 49.000 69.100 ;
        RECT 42.300 68.200 42.700 68.300 ;
        RECT 36.200 66.900 37.800 67.100 ;
        RECT 36.600 66.800 37.800 66.900 ;
        RECT 39.400 67.100 40.200 67.200 ;
        RECT 41.500 67.100 41.800 68.200 ;
        RECT 46.300 67.700 46.700 67.800 ;
        RECT 47.800 67.700 48.200 68.800 ;
        RECT 50.200 67.800 50.600 68.600 ;
        RECT 46.300 67.400 48.200 67.700 ;
        RECT 44.300 67.100 44.700 67.200 ;
        RECT 39.400 66.800 44.900 67.100 ;
        RECT 31.700 65.400 33.800 65.700 ;
        RECT 30.200 64.900 31.400 65.200 ;
        RECT 29.900 64.500 30.300 64.600 ;
        RECT 29.200 64.200 30.300 64.500 ;
        RECT 31.100 64.400 31.400 64.900 ;
        RECT 31.100 64.000 31.800 64.400 ;
        RECT 27.900 63.700 28.300 63.800 ;
        RECT 29.300 63.700 29.700 63.800 ;
        RECT 26.200 63.100 26.600 63.500 ;
        RECT 27.900 63.400 29.700 63.700 ;
        RECT 29.000 63.100 29.300 63.400 ;
        RECT 31.000 63.100 31.400 63.500 ;
        RECT 26.200 62.800 27.200 63.100 ;
        RECT 26.800 61.100 27.200 62.800 ;
        RECT 29.000 61.100 29.400 63.100 ;
        RECT 31.100 61.100 31.700 63.100 ;
        RECT 33.400 61.100 33.800 65.400 ;
        RECT 34.200 65.100 34.600 65.200 ;
        RECT 35.200 65.100 35.500 66.800 ;
        RECT 35.800 66.100 36.200 66.600 ;
        RECT 36.600 66.100 37.000 66.200 ;
        RECT 35.800 65.800 37.000 66.100 ;
        RECT 34.200 64.800 34.900 65.100 ;
        RECT 35.200 64.800 35.700 65.100 ;
        RECT 34.600 64.200 34.900 64.800 ;
        RECT 34.600 63.800 35.000 64.200 ;
        RECT 35.300 61.100 35.700 64.800 ;
        RECT 37.400 61.100 37.800 66.800 ;
        RECT 40.900 66.700 41.300 66.800 ;
        RECT 40.100 66.200 40.500 66.300 ;
        RECT 40.100 65.900 42.600 66.200 ;
        RECT 42.200 65.800 42.600 65.900 ;
        RECT 39.000 65.500 41.800 65.600 ;
        RECT 39.000 65.400 41.900 65.500 ;
        RECT 39.000 65.300 43.900 65.400 ;
        RECT 39.000 61.100 39.400 65.300 ;
        RECT 41.500 65.100 43.900 65.300 ;
        RECT 40.600 64.500 43.300 64.800 ;
        RECT 40.600 64.400 41.000 64.500 ;
        RECT 42.900 64.400 43.300 64.500 ;
        RECT 43.600 64.500 43.900 65.100 ;
        RECT 44.600 65.200 44.900 66.800 ;
        RECT 45.400 66.400 45.800 66.500 ;
        RECT 45.400 66.100 47.300 66.400 ;
        RECT 46.900 66.000 47.300 66.100 ;
        RECT 46.100 65.700 46.500 65.800 ;
        RECT 47.800 65.700 48.200 67.400 ;
        RECT 46.100 65.400 48.200 65.700 ;
        RECT 44.600 64.900 45.800 65.200 ;
        RECT 44.300 64.500 44.700 64.600 ;
        RECT 43.600 64.200 44.700 64.500 ;
        RECT 45.500 64.400 45.800 64.900 ;
        RECT 45.500 64.000 46.200 64.400 ;
        RECT 42.300 63.700 42.700 63.800 ;
        RECT 43.700 63.700 44.100 63.800 ;
        RECT 40.600 63.100 41.000 63.500 ;
        RECT 42.300 63.400 44.100 63.700 ;
        RECT 43.400 63.100 43.700 63.400 ;
        RECT 45.400 63.100 45.800 63.500 ;
        RECT 40.600 62.800 41.600 63.100 ;
        RECT 41.200 61.100 41.600 62.800 ;
        RECT 43.400 61.100 43.800 63.100 ;
        RECT 45.500 61.100 46.100 63.100 ;
        RECT 47.800 62.100 48.200 65.400 ;
        RECT 51.000 65.100 51.400 69.900 ;
        RECT 52.100 68.200 52.500 69.900 ;
        RECT 52.100 67.900 53.000 68.200 ;
        RECT 51.800 65.100 52.200 65.200 ;
        RECT 51.000 64.800 52.200 65.100 ;
        RECT 48.600 62.100 49.000 62.200 ;
        RECT 47.800 61.800 49.000 62.100 ;
        RECT 47.800 61.100 48.200 61.800 ;
        RECT 51.000 61.100 51.400 64.800 ;
        RECT 51.800 64.400 52.200 64.800 ;
        RECT 52.600 65.100 53.000 67.900 ;
        RECT 55.800 67.900 56.200 69.900 ;
        RECT 56.500 68.200 56.900 68.600 ;
        RECT 56.600 68.100 57.000 68.200 ;
        RECT 57.400 68.100 57.800 69.900 ;
        RECT 53.400 66.800 53.800 67.600 ;
        RECT 55.000 66.400 55.400 67.200 ;
        RECT 53.400 65.800 53.800 66.200 ;
        RECT 54.200 66.100 54.600 66.200 ;
        RECT 55.800 66.100 56.100 67.900 ;
        RECT 56.600 67.800 57.800 68.100 ;
        RECT 58.200 68.000 58.600 69.900 ;
        RECT 59.800 68.000 60.200 69.900 ;
        RECT 58.200 67.900 60.200 68.000 ;
        RECT 61.400 68.900 61.800 69.900 ;
        RECT 57.500 67.200 57.800 67.800 ;
        RECT 58.300 67.700 60.100 67.900 ;
        RECT 59.400 67.200 59.800 67.400 ;
        RECT 61.400 67.200 61.700 68.900 ;
        RECT 62.200 67.800 62.600 68.600 ;
        RECT 63.000 67.700 63.400 69.900 ;
        RECT 65.100 69.200 65.700 69.900 ;
        RECT 65.100 68.900 65.800 69.200 ;
        RECT 67.400 68.900 67.800 69.900 ;
        RECT 69.600 69.200 70.000 69.900 ;
        RECT 69.600 68.900 70.600 69.200 ;
        RECT 65.400 68.500 65.800 68.900 ;
        RECT 67.500 68.600 67.800 68.900 ;
        RECT 67.500 68.300 68.900 68.600 ;
        RECT 68.500 68.200 68.900 68.300 ;
        RECT 69.400 68.200 69.800 68.600 ;
        RECT 70.200 68.500 70.600 68.900 ;
        RECT 64.500 67.700 64.900 67.800 ;
        RECT 63.000 67.400 64.900 67.700 ;
        RECT 56.600 66.800 57.000 67.200 ;
        RECT 57.400 66.800 58.700 67.200 ;
        RECT 59.400 66.900 60.200 67.200 ;
        RECT 59.800 66.800 60.200 66.900 ;
        RECT 61.400 66.800 61.800 67.200 ;
        RECT 56.600 66.200 56.900 66.800 ;
        RECT 56.600 66.100 57.000 66.200 ;
        RECT 54.200 65.800 55.000 66.100 ;
        RECT 55.800 65.800 57.000 66.100 ;
        RECT 53.400 65.100 53.700 65.800 ;
        RECT 54.600 65.600 55.000 65.800 ;
        RECT 56.600 65.100 56.900 65.800 ;
        RECT 57.400 65.100 57.800 65.200 ;
        RECT 58.400 65.100 58.700 66.800 ;
        RECT 59.000 65.800 59.400 66.600 ;
        RECT 60.600 65.400 61.000 66.200 ;
        RECT 61.400 65.100 61.700 66.800 ;
        RECT 63.000 65.700 63.400 67.400 ;
        RECT 66.500 67.100 66.900 67.200 ;
        RECT 69.400 67.100 69.700 68.200 ;
        RECT 71.800 67.500 72.200 69.900 ;
        RECT 72.600 68.500 73.000 69.500 ;
        RECT 72.600 67.400 72.900 68.500 ;
        RECT 74.700 68.000 75.100 69.500 ;
        RECT 74.700 67.700 75.500 68.000 ;
        RECT 75.100 67.500 75.500 67.700 ;
        RECT 71.000 67.100 71.800 67.200 ;
        RECT 72.600 67.100 74.700 67.400 ;
        RECT 66.300 66.800 71.800 67.100 ;
        RECT 74.200 66.900 74.700 67.100 ;
        RECT 75.200 67.200 75.500 67.500 ;
        RECT 77.400 67.700 77.800 69.900 ;
        RECT 79.500 69.200 80.100 69.900 ;
        RECT 79.500 68.900 80.200 69.200 ;
        RECT 81.800 68.900 82.200 69.900 ;
        RECT 84.000 69.200 84.400 69.900 ;
        RECT 84.000 68.900 85.000 69.200 ;
        RECT 79.800 68.500 80.200 68.900 ;
        RECT 81.900 68.600 82.200 68.900 ;
        RECT 81.900 68.300 83.300 68.600 ;
        RECT 82.900 68.200 83.300 68.300 ;
        RECT 83.800 67.800 84.200 68.600 ;
        RECT 84.600 68.500 85.000 68.900 ;
        RECT 78.900 67.700 79.300 67.800 ;
        RECT 77.400 67.400 79.300 67.700 ;
        RECT 65.400 66.400 65.800 66.500 ;
        RECT 63.900 66.100 65.800 66.400 ;
        RECT 63.900 66.000 64.300 66.100 ;
        RECT 64.700 65.700 65.100 65.800 ;
        RECT 63.000 65.400 65.100 65.700 ;
        RECT 52.600 64.800 53.700 65.100 ;
        RECT 54.200 64.800 56.200 65.100 ;
        RECT 52.600 61.100 53.000 64.800 ;
        RECT 54.200 61.100 54.600 64.800 ;
        RECT 55.800 61.100 56.200 64.800 ;
        RECT 56.600 61.100 57.000 65.100 ;
        RECT 57.400 64.800 58.100 65.100 ;
        RECT 58.400 64.800 58.900 65.100 ;
        RECT 57.800 64.200 58.100 64.800 ;
        RECT 57.800 63.800 58.200 64.200 ;
        RECT 58.500 61.100 58.900 64.800 ;
        RECT 60.900 64.700 61.800 65.100 ;
        RECT 60.900 62.200 61.300 64.700 ;
        RECT 60.600 61.800 61.300 62.200 ;
        RECT 60.900 61.100 61.300 61.800 ;
        RECT 63.000 61.100 63.400 65.400 ;
        RECT 66.300 65.200 66.600 66.800 ;
        RECT 69.900 66.700 70.300 66.800 ;
        RECT 69.400 66.200 69.800 66.300 ;
        RECT 70.700 66.200 71.100 66.300 ;
        RECT 68.600 65.900 71.100 66.200 ;
        RECT 68.600 65.800 69.000 65.900 ;
        RECT 72.600 65.800 73.000 66.600 ;
        RECT 73.400 65.800 73.800 66.600 ;
        RECT 74.200 66.500 74.900 66.900 ;
        RECT 75.200 66.800 76.200 67.200 ;
        RECT 69.400 65.500 72.200 65.600 ;
        RECT 74.200 65.500 74.500 66.500 ;
        RECT 69.300 65.400 72.200 65.500 ;
        RECT 65.400 64.900 66.600 65.200 ;
        RECT 67.300 65.300 72.200 65.400 ;
        RECT 67.300 65.100 69.700 65.300 ;
        RECT 65.400 64.400 65.700 64.900 ;
        RECT 65.000 64.000 65.700 64.400 ;
        RECT 66.500 64.500 66.900 64.600 ;
        RECT 67.300 64.500 67.600 65.100 ;
        RECT 66.500 64.200 67.600 64.500 ;
        RECT 67.900 64.500 70.600 64.800 ;
        RECT 67.900 64.400 68.300 64.500 ;
        RECT 70.200 64.400 70.600 64.500 ;
        RECT 67.100 63.700 67.500 63.800 ;
        RECT 68.500 63.700 68.900 63.800 ;
        RECT 65.400 63.100 65.800 63.500 ;
        RECT 67.100 63.400 68.900 63.700 ;
        RECT 67.500 63.100 67.800 63.400 ;
        RECT 70.200 63.100 70.600 63.500 ;
        RECT 65.100 61.100 65.700 63.100 ;
        RECT 67.400 61.100 67.800 63.100 ;
        RECT 69.600 62.800 70.600 63.100 ;
        RECT 69.600 61.100 70.000 62.800 ;
        RECT 71.800 61.100 72.200 65.300 ;
        RECT 72.600 65.200 74.500 65.500 ;
        RECT 72.600 63.500 72.900 65.200 ;
        RECT 75.200 64.900 75.500 66.800 ;
        RECT 75.800 66.100 76.200 66.200 ;
        RECT 76.600 66.100 77.000 66.200 ;
        RECT 75.800 65.800 77.000 66.100 ;
        RECT 75.800 65.400 76.200 65.800 ;
        RECT 77.400 65.700 77.800 67.400 ;
        RECT 80.900 67.100 81.300 67.200 ;
        RECT 83.800 67.100 84.100 67.800 ;
        RECT 86.200 67.500 86.600 69.900 ;
        RECT 87.800 68.900 88.200 69.900 ;
        RECT 87.000 67.800 87.400 68.600 ;
        RECT 87.900 67.200 88.200 68.900 ;
        RECT 89.400 67.500 89.800 69.900 ;
        RECT 91.600 69.200 92.000 69.900 ;
        RECT 91.000 68.900 92.000 69.200 ;
        RECT 93.800 68.900 94.200 69.900 ;
        RECT 95.900 69.200 96.500 69.900 ;
        RECT 95.800 68.900 96.500 69.200 ;
        RECT 91.000 68.500 91.400 68.900 ;
        RECT 93.800 68.600 94.100 68.900 ;
        RECT 91.800 68.200 92.200 68.600 ;
        RECT 92.700 68.300 94.100 68.600 ;
        RECT 95.800 68.500 96.200 68.900 ;
        RECT 92.700 68.200 93.100 68.300 ;
        RECT 85.400 67.100 86.200 67.200 ;
        RECT 80.700 66.800 86.200 67.100 ;
        RECT 87.800 66.800 88.200 67.200 ;
        RECT 89.800 67.100 90.600 67.200 ;
        RECT 91.900 67.100 92.200 68.200 ;
        RECT 96.700 67.700 97.100 67.800 ;
        RECT 98.200 67.700 98.600 69.900 ;
        RECT 99.800 69.100 100.200 69.200 ;
        RECT 100.600 69.100 101.000 69.900 ;
        RECT 99.800 68.800 101.000 69.100 ;
        RECT 102.700 69.200 103.300 69.900 ;
        RECT 102.700 68.900 103.400 69.200 ;
        RECT 105.000 68.900 105.400 69.900 ;
        RECT 107.200 69.200 107.600 69.900 ;
        RECT 107.200 68.900 108.200 69.200 ;
        RECT 96.700 67.400 98.600 67.700 ;
        RECT 93.400 67.100 93.800 67.200 ;
        RECT 94.700 67.100 95.100 67.200 ;
        RECT 89.800 66.800 95.300 67.100 ;
        RECT 79.800 66.400 80.200 66.500 ;
        RECT 78.300 66.100 80.200 66.400 ;
        RECT 78.300 66.000 78.700 66.100 ;
        RECT 79.100 65.700 79.500 65.800 ;
        RECT 77.400 65.400 79.500 65.700 ;
        RECT 74.700 64.600 75.500 64.900 ;
        RECT 72.600 61.500 73.000 63.500 ;
        RECT 74.700 62.200 75.100 64.600 ;
        RECT 74.700 61.800 75.400 62.200 ;
        RECT 74.700 61.100 75.100 61.800 ;
        RECT 77.400 61.100 77.800 65.400 ;
        RECT 80.700 65.200 81.000 66.800 ;
        RECT 84.300 66.700 84.700 66.800 ;
        RECT 83.800 66.200 84.200 66.300 ;
        RECT 85.100 66.200 85.500 66.300 ;
        RECT 83.000 65.900 85.500 66.200 ;
        RECT 87.000 66.100 87.400 66.200 ;
        RECT 87.900 66.100 88.200 66.800 ;
        RECT 91.300 66.700 91.700 66.800 ;
        RECT 90.500 66.200 90.900 66.300 ;
        RECT 91.800 66.200 92.200 66.300 ;
        RECT 83.000 65.800 83.400 65.900 ;
        RECT 87.000 65.800 88.200 66.100 ;
        RECT 83.800 65.500 86.600 65.600 ;
        RECT 83.700 65.400 86.600 65.500 ;
        RECT 79.800 64.900 81.000 65.200 ;
        RECT 81.700 65.300 86.600 65.400 ;
        RECT 81.700 65.100 84.100 65.300 ;
        RECT 79.800 64.400 80.100 64.900 ;
        RECT 79.400 64.000 80.100 64.400 ;
        RECT 80.900 64.500 81.300 64.600 ;
        RECT 81.700 64.500 82.000 65.100 ;
        RECT 80.900 64.200 82.000 64.500 ;
        RECT 82.300 64.500 85.000 64.800 ;
        RECT 82.300 64.400 82.700 64.500 ;
        RECT 84.600 64.400 85.000 64.500 ;
        RECT 81.500 63.700 81.900 63.800 ;
        RECT 82.900 63.700 83.300 63.800 ;
        RECT 79.800 63.100 80.200 63.500 ;
        RECT 81.500 63.400 83.300 63.700 ;
        RECT 81.900 63.100 82.200 63.400 ;
        RECT 84.600 63.100 85.000 63.500 ;
        RECT 79.500 61.100 80.100 63.100 ;
        RECT 81.800 61.100 82.200 63.100 ;
        RECT 84.000 62.800 85.000 63.100 ;
        RECT 84.000 61.100 84.400 62.800 ;
        RECT 86.200 61.100 86.600 65.300 ;
        RECT 87.900 65.100 88.200 65.800 ;
        RECT 88.600 65.400 89.000 66.200 ;
        RECT 90.500 65.900 93.000 66.200 ;
        RECT 92.600 65.800 93.000 65.900 ;
        RECT 89.400 65.500 92.200 65.600 ;
        RECT 89.400 65.400 92.300 65.500 ;
        RECT 89.400 65.300 94.300 65.400 ;
        RECT 87.800 64.700 88.700 65.100 ;
        RECT 88.300 61.100 88.700 64.700 ;
        RECT 89.400 61.100 89.800 65.300 ;
        RECT 91.900 65.100 94.300 65.300 ;
        RECT 91.000 64.500 93.700 64.800 ;
        RECT 91.000 64.400 91.400 64.500 ;
        RECT 93.300 64.400 93.700 64.500 ;
        RECT 94.000 64.500 94.300 65.100 ;
        RECT 95.000 65.200 95.300 66.800 ;
        RECT 95.800 66.400 96.200 66.500 ;
        RECT 95.800 66.100 97.700 66.400 ;
        RECT 97.300 66.000 97.700 66.100 ;
        RECT 96.500 65.700 96.900 65.800 ;
        RECT 98.200 65.700 98.600 67.400 ;
        RECT 96.500 65.400 98.600 65.700 ;
        RECT 95.000 64.900 96.200 65.200 ;
        RECT 94.700 64.500 95.100 64.600 ;
        RECT 94.000 64.200 95.100 64.500 ;
        RECT 95.900 64.400 96.200 64.900 ;
        RECT 95.900 64.000 96.600 64.400 ;
        RECT 92.700 63.700 93.100 63.800 ;
        RECT 94.100 63.700 94.500 63.800 ;
        RECT 91.000 63.100 91.400 63.500 ;
        RECT 92.700 63.400 94.500 63.700 ;
        RECT 93.800 63.100 94.100 63.400 ;
        RECT 95.800 63.100 96.200 63.500 ;
        RECT 91.000 62.800 92.000 63.100 ;
        RECT 91.600 61.100 92.000 62.800 ;
        RECT 93.800 61.100 94.200 63.100 ;
        RECT 95.900 61.100 96.500 63.100 ;
        RECT 98.200 61.100 98.600 65.400 ;
        RECT 100.600 67.700 101.000 68.800 ;
        RECT 103.000 68.500 103.400 68.900 ;
        RECT 105.100 68.600 105.400 68.900 ;
        RECT 105.100 68.300 106.500 68.600 ;
        RECT 106.100 68.200 106.500 68.300 ;
        RECT 103.800 67.800 104.200 68.200 ;
        RECT 107.000 67.800 107.400 68.600 ;
        RECT 107.800 68.500 108.200 68.900 ;
        RECT 102.100 67.700 102.500 67.800 ;
        RECT 100.600 67.400 102.500 67.700 ;
        RECT 100.600 65.700 101.000 67.400 ;
        RECT 103.800 67.200 104.100 67.800 ;
        RECT 103.800 67.100 104.500 67.200 ;
        RECT 107.000 67.100 107.300 67.800 ;
        RECT 109.400 67.500 109.800 69.900 ;
        RECT 110.200 67.800 110.600 68.600 ;
        RECT 111.000 68.100 111.400 69.900 ;
        RECT 112.600 68.900 113.000 69.900 ;
        RECT 111.800 68.100 112.200 68.600 ;
        RECT 111.000 67.800 112.200 68.100 ;
        RECT 108.600 67.100 109.400 67.200 ;
        RECT 103.800 66.800 109.400 67.100 ;
        RECT 103.000 66.400 103.400 66.500 ;
        RECT 101.500 66.100 103.400 66.400 ;
        RECT 101.500 66.000 101.900 66.100 ;
        RECT 102.300 65.700 102.700 65.800 ;
        RECT 100.600 65.400 102.700 65.700 ;
        RECT 100.600 61.100 101.000 65.400 ;
        RECT 103.900 65.200 104.200 66.800 ;
        RECT 107.500 66.700 107.900 66.800 ;
        RECT 107.000 66.200 107.400 66.300 ;
        RECT 108.300 66.200 108.700 66.300 ;
        RECT 106.200 65.900 108.700 66.200 ;
        RECT 106.200 65.800 106.600 65.900 ;
        RECT 107.000 65.500 109.800 65.600 ;
        RECT 106.900 65.400 109.800 65.500 ;
        RECT 103.000 64.900 104.200 65.200 ;
        RECT 104.900 65.300 109.800 65.400 ;
        RECT 104.900 65.100 107.300 65.300 ;
        RECT 103.000 64.400 103.300 64.900 ;
        RECT 102.600 64.000 103.300 64.400 ;
        RECT 104.100 64.500 104.500 64.600 ;
        RECT 104.900 64.500 105.200 65.100 ;
        RECT 104.100 64.200 105.200 64.500 ;
        RECT 105.500 64.500 108.200 64.800 ;
        RECT 105.500 64.400 105.900 64.500 ;
        RECT 107.800 64.400 108.200 64.500 ;
        RECT 104.700 63.700 105.100 63.800 ;
        RECT 106.100 63.700 106.500 63.800 ;
        RECT 103.000 63.100 103.400 63.500 ;
        RECT 104.700 63.400 106.500 63.700 ;
        RECT 105.100 63.100 105.400 63.400 ;
        RECT 107.800 63.100 108.200 63.500 ;
        RECT 102.700 61.100 103.300 63.100 ;
        RECT 105.000 61.100 105.400 63.100 ;
        RECT 107.200 62.800 108.200 63.100 ;
        RECT 107.200 61.100 107.600 62.800 ;
        RECT 109.400 61.100 109.800 65.300 ;
        RECT 111.000 61.100 111.400 67.800 ;
        RECT 112.700 67.200 113.000 68.900 ;
        RECT 114.200 67.500 114.600 69.900 ;
        RECT 116.400 69.200 116.800 69.900 ;
        RECT 115.800 68.900 116.800 69.200 ;
        RECT 118.600 68.900 119.000 69.900 ;
        RECT 120.700 69.200 121.300 69.900 ;
        RECT 120.600 68.900 121.300 69.200 ;
        RECT 115.800 68.500 116.200 68.900 ;
        RECT 118.600 68.600 118.900 68.900 ;
        RECT 116.600 67.800 117.000 68.600 ;
        RECT 117.500 68.300 118.900 68.600 ;
        RECT 120.600 68.500 121.000 68.900 ;
        RECT 117.500 68.200 117.900 68.300 ;
        RECT 112.600 66.800 113.000 67.200 ;
        RECT 114.600 67.100 115.400 67.200 ;
        RECT 116.700 67.100 117.000 67.800 ;
        RECT 121.500 67.700 121.900 67.800 ;
        RECT 123.000 67.700 123.400 69.900 ;
        RECT 121.500 67.400 123.400 67.700 ;
        RECT 119.500 67.100 119.900 67.200 ;
        RECT 114.600 66.800 120.100 67.100 ;
        RECT 112.700 65.100 113.000 66.800 ;
        RECT 116.100 66.700 116.500 66.800 ;
        RECT 115.300 66.200 115.700 66.300 ;
        RECT 113.400 65.400 113.800 66.200 ;
        RECT 115.300 66.100 117.800 66.200 ;
        RECT 119.000 66.100 119.400 66.200 ;
        RECT 115.300 65.900 119.400 66.100 ;
        RECT 117.400 65.800 119.400 65.900 ;
        RECT 114.200 65.500 117.000 65.600 ;
        RECT 114.200 65.400 117.100 65.500 ;
        RECT 114.200 65.300 119.100 65.400 ;
        RECT 112.600 64.700 113.500 65.100 ;
        RECT 113.100 61.100 113.500 64.700 ;
        RECT 114.200 61.100 114.600 65.300 ;
        RECT 116.700 65.100 119.100 65.300 ;
        RECT 115.800 64.500 118.500 64.800 ;
        RECT 115.800 64.400 116.200 64.500 ;
        RECT 118.100 64.400 118.500 64.500 ;
        RECT 118.800 64.500 119.100 65.100 ;
        RECT 119.800 65.200 120.100 66.800 ;
        RECT 120.600 66.400 121.000 66.500 ;
        RECT 120.600 66.100 122.500 66.400 ;
        RECT 122.100 66.000 122.500 66.100 ;
        RECT 121.300 65.700 121.700 65.800 ;
        RECT 123.000 65.700 123.400 67.400 ;
        RECT 124.600 67.600 125.000 69.900 ;
        RECT 126.200 67.600 126.600 69.900 ;
        RECT 127.800 67.600 128.200 69.900 ;
        RECT 129.400 67.600 129.800 69.900 ;
        RECT 124.600 67.200 125.500 67.600 ;
        RECT 126.200 67.200 127.300 67.600 ;
        RECT 127.800 67.200 128.900 67.600 ;
        RECT 129.400 67.200 130.600 67.600 ;
        RECT 131.000 67.500 131.400 69.900 ;
        RECT 133.200 69.200 133.600 69.900 ;
        RECT 132.600 68.900 133.600 69.200 ;
        RECT 135.400 68.900 135.800 69.900 ;
        RECT 137.500 69.200 138.100 69.900 ;
        RECT 137.400 68.900 138.100 69.200 ;
        RECT 132.600 68.500 133.000 68.900 ;
        RECT 135.400 68.600 135.700 68.900 ;
        RECT 133.400 67.800 133.800 68.600 ;
        RECT 134.300 68.300 135.700 68.600 ;
        RECT 137.400 68.500 137.800 68.900 ;
        RECT 134.300 68.200 134.700 68.300 ;
        RECT 125.100 66.900 125.500 67.200 ;
        RECT 126.900 66.900 127.300 67.200 ;
        RECT 128.500 66.900 128.900 67.200 ;
        RECT 125.100 66.500 126.400 66.900 ;
        RECT 126.900 66.500 128.100 66.900 ;
        RECT 128.500 66.500 129.800 66.900 ;
        RECT 125.100 65.800 125.500 66.500 ;
        RECT 126.900 65.800 127.300 66.500 ;
        RECT 128.500 65.800 128.900 66.500 ;
        RECT 130.200 65.800 130.600 67.200 ;
        RECT 131.400 67.100 132.200 67.200 ;
        RECT 133.500 67.100 133.800 67.800 ;
        RECT 138.300 67.700 138.700 67.800 ;
        RECT 139.800 67.700 140.200 69.900 ;
        RECT 138.300 67.400 140.200 67.700 ;
        RECT 136.300 67.100 136.700 67.200 ;
        RECT 131.400 66.800 136.900 67.100 ;
        RECT 132.900 66.700 133.300 66.800 ;
        RECT 132.100 66.200 132.500 66.300 ;
        RECT 132.100 65.900 134.600 66.200 ;
        RECT 134.200 65.800 134.600 65.900 ;
        RECT 121.300 65.400 123.400 65.700 ;
        RECT 119.800 64.900 121.000 65.200 ;
        RECT 119.500 64.500 119.900 64.600 ;
        RECT 118.800 64.200 119.900 64.500 ;
        RECT 120.700 64.400 121.000 64.900 ;
        RECT 120.700 64.000 121.400 64.400 ;
        RECT 117.500 63.700 117.900 63.800 ;
        RECT 118.900 63.700 119.300 63.800 ;
        RECT 115.800 63.100 116.200 63.500 ;
        RECT 117.500 63.400 119.300 63.700 ;
        RECT 118.600 63.100 118.900 63.400 ;
        RECT 120.600 63.100 121.000 63.500 ;
        RECT 115.800 62.800 116.800 63.100 ;
        RECT 116.400 61.100 116.800 62.800 ;
        RECT 118.600 61.100 119.000 63.100 ;
        RECT 120.700 61.100 121.300 63.100 ;
        RECT 123.000 61.100 123.400 65.400 ;
        RECT 124.600 65.400 125.500 65.800 ;
        RECT 126.200 65.400 127.300 65.800 ;
        RECT 127.800 65.400 128.900 65.800 ;
        RECT 129.400 65.400 130.600 65.800 ;
        RECT 131.000 65.500 133.800 65.600 ;
        RECT 131.000 65.400 133.900 65.500 ;
        RECT 124.600 61.100 125.000 65.400 ;
        RECT 126.200 61.100 126.600 65.400 ;
        RECT 127.800 61.100 128.200 65.400 ;
        RECT 129.400 61.100 129.800 65.400 ;
        RECT 131.000 65.300 135.900 65.400 ;
        RECT 131.000 61.100 131.400 65.300 ;
        RECT 133.500 65.100 135.900 65.300 ;
        RECT 132.600 64.500 135.300 64.800 ;
        RECT 132.600 64.400 133.000 64.500 ;
        RECT 134.900 64.400 135.300 64.500 ;
        RECT 135.600 64.500 135.900 65.100 ;
        RECT 136.600 65.200 136.900 66.800 ;
        RECT 137.400 66.400 137.800 66.500 ;
        RECT 137.400 66.100 139.300 66.400 ;
        RECT 138.900 66.000 139.300 66.100 ;
        RECT 138.100 65.700 138.500 65.800 ;
        RECT 139.800 65.700 140.200 67.400 ;
        RECT 141.400 67.600 141.800 69.900 ;
        RECT 143.000 67.600 143.400 69.900 ;
        RECT 144.600 67.600 145.000 69.900 ;
        RECT 146.200 67.600 146.600 69.900 ;
        RECT 141.400 67.200 142.300 67.600 ;
        RECT 143.000 67.200 144.100 67.600 ;
        RECT 144.600 67.200 145.700 67.600 ;
        RECT 146.200 67.200 147.400 67.600 ;
        RECT 141.900 66.900 142.300 67.200 ;
        RECT 143.700 66.900 144.100 67.200 ;
        RECT 145.300 66.900 145.700 67.200 ;
        RECT 141.900 66.500 143.200 66.900 ;
        RECT 143.700 66.500 144.900 66.900 ;
        RECT 145.300 66.500 146.600 66.900 ;
        RECT 141.900 65.800 142.300 66.500 ;
        RECT 143.700 65.800 144.100 66.500 ;
        RECT 145.300 65.800 145.700 66.500 ;
        RECT 147.000 65.800 147.400 67.200 ;
        RECT 138.100 65.400 140.200 65.700 ;
        RECT 136.600 64.900 137.800 65.200 ;
        RECT 136.300 64.500 136.700 64.600 ;
        RECT 135.600 64.200 136.700 64.500 ;
        RECT 137.500 64.400 137.800 64.900 ;
        RECT 137.500 64.000 138.200 64.400 ;
        RECT 134.300 63.700 134.700 63.800 ;
        RECT 135.700 63.700 136.100 63.800 ;
        RECT 132.600 63.100 133.000 63.500 ;
        RECT 134.300 63.400 136.100 63.700 ;
        RECT 135.400 63.100 135.700 63.400 ;
        RECT 137.400 63.100 137.800 63.500 ;
        RECT 132.600 62.800 133.600 63.100 ;
        RECT 133.200 61.100 133.600 62.800 ;
        RECT 135.400 61.100 135.800 63.100 ;
        RECT 137.500 61.100 138.100 63.100 ;
        RECT 139.800 61.100 140.200 65.400 ;
        RECT 141.400 65.400 142.300 65.800 ;
        RECT 143.000 65.400 144.100 65.800 ;
        RECT 144.600 65.400 145.700 65.800 ;
        RECT 146.200 65.400 147.400 65.800 ;
        RECT 149.400 66.200 149.800 69.900 ;
        RECT 151.000 67.600 151.400 69.900 ;
        RECT 152.100 68.400 152.500 69.900 ;
        RECT 150.300 67.300 151.400 67.600 ;
        RECT 151.800 67.900 152.500 68.400 ;
        RECT 154.200 67.900 154.600 69.900 ;
        RECT 141.400 61.100 141.800 65.400 ;
        RECT 143.000 61.100 143.400 65.400 ;
        RECT 144.600 61.100 145.000 65.400 ;
        RECT 146.200 61.100 146.600 65.400 ;
        RECT 149.400 65.100 149.700 66.200 ;
        RECT 150.300 65.800 150.600 67.300 ;
        RECT 151.000 66.100 151.400 66.600 ;
        RECT 151.800 66.200 152.100 67.900 ;
        RECT 154.200 67.800 154.500 67.900 ;
        RECT 153.600 67.600 154.500 67.800 ;
        RECT 152.400 67.500 154.500 67.600 ;
        RECT 155.000 67.600 155.400 69.900 ;
        RECT 152.400 67.300 153.900 67.500 ;
        RECT 155.000 67.300 156.100 67.600 ;
        RECT 152.400 67.200 152.800 67.300 ;
        RECT 151.800 66.100 152.200 66.200 ;
        RECT 151.000 65.800 152.200 66.100 ;
        RECT 150.000 65.400 150.600 65.800 ;
        RECT 150.300 65.100 150.600 65.400 ;
        RECT 151.800 65.100 152.100 65.800 ;
        RECT 152.500 65.500 152.800 67.200 ;
        RECT 153.200 66.900 153.600 67.000 ;
        RECT 153.200 66.600 153.700 66.900 ;
        RECT 153.400 66.200 153.700 66.600 ;
        RECT 154.200 66.400 154.600 67.200 ;
        RECT 153.400 65.800 153.800 66.200 ;
        RECT 155.000 65.800 155.400 66.600 ;
        RECT 155.800 65.800 156.100 67.300 ;
        RECT 156.600 66.200 157.000 69.900 ;
        RECT 157.700 68.400 158.100 69.900 ;
        RECT 152.500 65.200 153.700 65.500 ;
        RECT 149.400 61.100 149.800 65.100 ;
        RECT 150.300 64.800 151.400 65.100 ;
        RECT 151.000 61.100 151.400 64.800 ;
        RECT 151.800 61.100 152.200 65.100 ;
        RECT 153.400 63.100 153.700 65.200 ;
        RECT 155.800 65.400 156.400 65.800 ;
        RECT 155.800 65.100 156.100 65.400 ;
        RECT 156.700 65.100 157.000 66.200 ;
        RECT 155.000 64.800 156.100 65.100 ;
        RECT 153.400 61.100 153.800 63.100 ;
        RECT 155.000 61.100 155.400 64.800 ;
        RECT 156.600 61.100 157.000 65.100 ;
        RECT 157.400 67.900 158.100 68.400 ;
        RECT 159.800 67.900 160.200 69.900 ;
        RECT 160.900 68.200 161.300 69.900 ;
        RECT 163.600 69.200 164.000 69.900 ;
        RECT 163.600 68.800 164.200 69.200 ;
        RECT 157.400 66.200 157.700 67.900 ;
        RECT 159.800 67.800 160.100 67.900 ;
        RECT 159.200 67.600 160.100 67.800 ;
        RECT 158.000 67.500 160.100 67.600 ;
        RECT 160.600 67.800 161.800 68.200 ;
        RECT 158.000 67.300 159.500 67.500 ;
        RECT 158.000 67.200 158.400 67.300 ;
        RECT 160.600 67.200 160.900 67.800 ;
        RECT 157.400 65.800 157.800 66.200 ;
        RECT 157.400 65.100 157.700 65.800 ;
        RECT 158.100 65.500 158.400 67.200 ;
        RECT 158.800 66.900 159.200 67.000 ;
        RECT 158.800 66.600 159.300 66.900 ;
        RECT 159.000 66.200 159.300 66.600 ;
        RECT 159.800 66.400 160.200 67.200 ;
        RECT 160.600 66.800 161.000 67.200 ;
        RECT 159.000 65.800 159.400 66.200 ;
        RECT 158.100 65.200 159.300 65.500 ;
        RECT 157.400 61.100 157.800 65.100 ;
        RECT 159.000 63.100 159.300 65.200 ;
        RECT 160.600 64.400 161.000 65.200 ;
        RECT 159.000 61.100 159.400 63.100 ;
        RECT 161.400 61.100 161.800 67.800 ;
        RECT 162.200 66.800 162.600 67.600 ;
        RECT 163.600 67.100 164.000 68.800 ;
        RECT 163.100 66.900 164.000 67.100 ;
        RECT 163.100 66.800 163.900 66.900 ;
        RECT 166.200 66.800 166.600 67.600 ;
        RECT 167.000 67.100 167.400 69.900 ;
        RECT 169.100 68.200 169.500 69.900 ;
        RECT 168.600 67.800 169.700 68.200 ;
        RECT 167.800 67.100 168.200 67.600 ;
        RECT 167.000 66.800 168.200 67.100 ;
        RECT 163.100 65.200 163.400 66.800 ;
        RECT 164.200 65.800 165.000 66.200 ;
        RECT 167.000 66.100 167.400 66.800 ;
        RECT 165.400 65.800 167.400 66.100 ;
        RECT 163.000 64.800 163.400 65.200 ;
        RECT 165.400 64.800 165.800 65.800 ;
        RECT 163.100 63.500 163.400 64.800 ;
        RECT 163.800 63.800 164.200 64.600 ;
        RECT 163.100 63.200 164.900 63.500 ;
        RECT 163.100 63.100 163.400 63.200 ;
        RECT 163.000 61.100 163.400 63.100 ;
        RECT 164.600 63.100 164.900 63.200 ;
        RECT 164.600 61.100 165.000 63.100 ;
        RECT 167.000 61.100 167.400 65.800 ;
        RECT 168.600 61.100 169.000 67.800 ;
        RECT 169.400 67.200 169.700 67.800 ;
        RECT 171.000 68.100 171.400 69.900 ;
        RECT 172.600 68.900 173.000 69.900 ;
        RECT 171.800 68.100 172.200 68.200 ;
        RECT 171.000 67.800 172.200 68.100 ;
        RECT 169.400 66.800 169.800 67.200 ;
        RECT 170.200 66.800 170.600 67.600 ;
        RECT 171.000 66.100 171.400 67.800 ;
        RECT 172.600 67.200 172.900 68.900 ;
        RECT 173.400 67.800 173.800 68.600 ;
        RECT 174.200 67.900 174.600 69.900 ;
        RECT 175.000 68.000 175.400 69.900 ;
        RECT 176.600 68.000 177.000 69.900 ;
        RECT 175.000 67.900 177.000 68.000 ;
        RECT 178.200 68.900 178.600 69.900 ;
        RECT 174.300 67.200 174.600 67.900 ;
        RECT 175.100 67.700 176.900 67.900 ;
        RECT 176.200 67.200 176.600 67.400 ;
        RECT 178.200 67.200 178.500 68.900 ;
        RECT 179.000 67.800 179.400 68.600 ;
        RECT 179.800 67.500 180.200 69.900 ;
        RECT 182.000 69.200 182.400 69.900 ;
        RECT 181.400 68.900 182.400 69.200 ;
        RECT 184.200 68.900 184.600 69.900 ;
        RECT 186.300 69.200 186.900 69.900 ;
        RECT 186.200 68.900 186.900 69.200 ;
        RECT 181.400 68.500 181.800 68.900 ;
        RECT 184.200 68.600 184.500 68.900 ;
        RECT 182.200 68.200 182.600 68.600 ;
        RECT 183.100 68.300 184.500 68.600 ;
        RECT 186.200 68.500 186.600 68.900 ;
        RECT 183.100 68.200 183.500 68.300 ;
        RECT 172.600 66.800 173.000 67.200 ;
        RECT 174.200 66.800 175.500 67.200 ;
        RECT 176.200 66.900 177.000 67.200 ;
        RECT 176.600 66.800 177.000 66.900 ;
        RECT 178.200 66.800 178.600 67.200 ;
        RECT 180.200 67.100 181.000 67.200 ;
        RECT 182.300 67.100 182.600 68.200 ;
        RECT 187.100 67.700 187.500 67.800 ;
        RECT 188.600 67.700 189.000 69.900 ;
        RECT 187.100 67.400 189.000 67.700 ;
        RECT 185.100 67.100 185.500 67.200 ;
        RECT 180.200 66.800 185.700 67.100 ;
        RECT 171.800 66.100 172.200 66.200 ;
        RECT 171.000 65.800 172.200 66.100 ;
        RECT 169.400 64.400 169.800 65.200 ;
        RECT 171.000 61.100 171.400 65.800 ;
        RECT 171.800 65.400 172.200 65.800 ;
        RECT 172.600 66.100 172.900 66.800 ;
        RECT 173.400 66.100 173.800 66.200 ;
        RECT 172.600 65.800 173.800 66.100 ;
        RECT 172.600 65.100 172.900 65.800 ;
        RECT 175.200 65.200 175.500 66.800 ;
        RECT 175.800 65.800 176.200 66.600 ;
        RECT 176.600 66.100 177.000 66.200 ;
        RECT 177.400 66.100 177.800 66.200 ;
        RECT 176.600 65.800 177.800 66.100 ;
        RECT 177.400 65.400 177.800 65.800 ;
        RECT 174.200 65.100 174.600 65.200 ;
        RECT 172.100 64.700 173.000 65.100 ;
        RECT 174.200 64.800 174.900 65.100 ;
        RECT 175.200 64.800 176.200 65.200 ;
        RECT 178.200 65.100 178.500 66.800 ;
        RECT 181.700 66.700 182.100 66.800 ;
        RECT 180.900 66.200 181.300 66.300 ;
        RECT 182.200 66.200 182.600 66.300 ;
        RECT 180.900 65.900 183.400 66.200 ;
        RECT 183.000 65.800 183.400 65.900 ;
        RECT 179.800 65.500 182.600 65.600 ;
        RECT 179.800 65.400 182.700 65.500 ;
        RECT 179.800 65.300 184.700 65.400 ;
        RECT 172.100 61.100 172.500 64.700 ;
        RECT 174.600 64.200 174.900 64.800 ;
        RECT 174.600 63.800 175.000 64.200 ;
        RECT 175.300 61.100 175.700 64.800 ;
        RECT 177.700 64.700 178.600 65.100 ;
        RECT 177.700 62.200 178.100 64.700 ;
        RECT 177.700 61.800 178.600 62.200 ;
        RECT 177.700 61.100 178.100 61.800 ;
        RECT 179.800 61.100 180.200 65.300 ;
        RECT 182.300 65.100 184.700 65.300 ;
        RECT 181.400 64.500 184.100 64.800 ;
        RECT 181.400 64.400 181.800 64.500 ;
        RECT 183.700 64.400 184.100 64.500 ;
        RECT 184.400 64.500 184.700 65.100 ;
        RECT 185.400 65.200 185.700 66.800 ;
        RECT 186.200 66.400 186.600 66.500 ;
        RECT 186.200 66.100 188.100 66.400 ;
        RECT 187.700 66.000 188.100 66.100 ;
        RECT 186.900 65.700 187.300 65.800 ;
        RECT 188.600 65.700 189.000 67.400 ;
        RECT 189.400 67.600 189.800 69.900 ;
        RECT 191.800 67.600 192.200 69.900 ;
        RECT 189.400 67.300 190.500 67.600 ;
        RECT 191.800 67.300 192.900 67.600 ;
        RECT 186.900 65.400 189.000 65.700 ;
        RECT 185.400 64.900 186.600 65.200 ;
        RECT 185.100 64.500 185.500 64.600 ;
        RECT 184.400 64.200 185.500 64.500 ;
        RECT 186.300 64.400 186.600 64.900 ;
        RECT 186.300 64.200 187.000 64.400 ;
        RECT 186.300 64.000 187.400 64.200 ;
        RECT 186.700 63.800 187.400 64.000 ;
        RECT 183.100 63.700 183.500 63.800 ;
        RECT 184.500 63.700 184.900 63.800 ;
        RECT 181.400 63.100 181.800 63.500 ;
        RECT 183.100 63.400 184.900 63.700 ;
        RECT 184.200 63.100 184.500 63.400 ;
        RECT 186.200 63.100 186.600 63.500 ;
        RECT 181.400 62.800 182.400 63.100 ;
        RECT 182.000 61.100 182.400 62.800 ;
        RECT 184.200 61.100 184.600 63.100 ;
        RECT 186.300 61.100 186.900 63.100 ;
        RECT 188.600 61.100 189.000 65.400 ;
        RECT 190.200 65.800 190.500 67.300 ;
        RECT 192.600 65.800 192.900 67.300 ;
        RECT 190.200 65.400 190.800 65.800 ;
        RECT 192.600 65.400 193.200 65.800 ;
        RECT 190.200 65.100 190.500 65.400 ;
        RECT 192.600 65.100 192.900 65.400 ;
        RECT 189.400 64.800 190.500 65.100 ;
        RECT 191.800 64.800 192.900 65.100 ;
        RECT 189.400 61.100 189.800 64.800 ;
        RECT 191.800 61.100 192.200 64.800 ;
        RECT 1.400 55.600 1.800 59.900 ;
        RECT 3.000 55.600 3.400 59.900 ;
        RECT 4.600 55.600 5.000 59.900 ;
        RECT 6.200 55.600 6.600 59.900 ;
        RECT 9.100 56.300 9.500 59.900 ;
        RECT 8.600 55.900 9.500 56.300 ;
        RECT 10.200 57.500 10.600 59.500 ;
        RECT 1.400 55.200 2.300 55.600 ;
        RECT 3.000 55.200 4.100 55.600 ;
        RECT 4.600 55.200 5.700 55.600 ;
        RECT 6.200 55.200 7.400 55.600 ;
        RECT 1.900 54.500 2.300 55.200 ;
        RECT 3.700 54.500 4.100 55.200 ;
        RECT 5.300 54.500 5.700 55.200 ;
        RECT 1.900 54.100 3.200 54.500 ;
        RECT 3.700 54.100 4.900 54.500 ;
        RECT 5.300 54.100 6.600 54.500 ;
        RECT 1.900 53.800 2.300 54.100 ;
        RECT 3.700 53.800 4.100 54.100 ;
        RECT 5.300 53.800 5.700 54.100 ;
        RECT 7.000 53.800 7.400 55.200 ;
        RECT 8.700 54.200 9.000 55.900 ;
        RECT 10.200 55.800 10.500 57.500 ;
        RECT 12.300 57.200 12.700 59.900 ;
        RECT 12.300 56.800 13.000 57.200 ;
        RECT 12.300 56.400 12.700 56.800 ;
        RECT 12.300 56.100 13.100 56.400 ;
        RECT 9.400 54.800 9.800 55.600 ;
        RECT 10.200 55.500 12.100 55.800 ;
        RECT 10.200 54.400 10.600 55.200 ;
        RECT 11.000 54.400 11.400 55.200 ;
        RECT 11.800 54.500 12.100 55.500 ;
        RECT 8.600 53.800 9.000 54.200 ;
        RECT 11.800 54.100 12.500 54.500 ;
        RECT 12.800 54.200 13.100 56.100 ;
        RECT 13.400 54.800 13.800 55.600 ;
        RECT 11.800 53.900 12.300 54.100 ;
        RECT 1.400 53.400 2.300 53.800 ;
        RECT 3.000 53.400 4.100 53.800 ;
        RECT 4.600 53.400 5.700 53.800 ;
        RECT 6.200 53.400 7.400 53.800 ;
        RECT 1.400 51.100 1.800 53.400 ;
        RECT 3.000 51.100 3.400 53.400 ;
        RECT 4.600 51.100 5.000 53.400 ;
        RECT 6.200 51.100 6.600 53.400 ;
        RECT 7.800 52.400 8.200 53.200 ;
        RECT 8.700 53.100 9.000 53.800 ;
        RECT 10.200 53.600 12.300 53.900 ;
        RECT 12.800 53.800 13.800 54.200 ;
        RECT 9.400 53.100 9.800 53.200 ;
        RECT 8.600 52.800 9.800 53.100 ;
        RECT 8.700 52.100 9.000 52.800 ;
        RECT 8.600 51.100 9.000 52.100 ;
        RECT 10.200 52.500 10.500 53.600 ;
        RECT 12.800 53.500 13.100 53.800 ;
        RECT 12.700 53.300 13.100 53.500 ;
        RECT 15.000 53.400 15.400 54.200 ;
        RECT 12.300 53.000 13.100 53.300 ;
        RECT 15.800 53.100 16.200 59.900 ;
        RECT 16.600 55.800 17.000 56.600 ;
        RECT 18.200 56.400 18.600 59.900 ;
        RECT 18.100 55.900 18.600 56.400 ;
        RECT 19.800 56.200 20.200 59.900 ;
        RECT 21.900 56.300 22.300 59.900 ;
        RECT 18.900 55.900 20.200 56.200 ;
        RECT 21.400 55.900 22.300 56.300 ;
        RECT 23.000 57.500 23.400 59.500 ;
        RECT 18.100 54.200 18.400 55.900 ;
        RECT 18.900 54.900 19.200 55.900 ;
        RECT 18.700 54.500 19.200 54.900 ;
        RECT 16.600 54.100 17.000 54.200 ;
        RECT 18.100 54.100 18.600 54.200 ;
        RECT 16.600 53.800 18.600 54.100 ;
        RECT 18.100 53.100 18.400 53.800 ;
        RECT 18.900 53.700 19.200 54.500 ;
        RECT 19.700 54.800 20.200 55.200 ;
        RECT 19.700 54.400 20.100 54.800 ;
        RECT 21.500 54.200 21.800 55.900 ;
        RECT 23.000 55.800 23.300 57.500 ;
        RECT 25.100 56.400 25.500 59.900 ;
        RECT 25.100 56.100 25.900 56.400 ;
        RECT 22.200 54.800 22.600 55.600 ;
        RECT 23.000 55.500 24.900 55.800 ;
        RECT 23.000 54.400 23.400 55.200 ;
        RECT 23.800 54.400 24.200 55.200 ;
        RECT 24.600 54.500 24.900 55.500 ;
        RECT 21.400 53.800 21.800 54.200 ;
        RECT 24.600 54.100 25.300 54.500 ;
        RECT 25.600 54.200 25.900 56.100 ;
        RECT 26.200 55.100 26.600 55.600 ;
        RECT 27.800 55.100 28.200 55.200 ;
        RECT 26.200 54.800 28.200 55.100 ;
        RECT 24.600 53.900 25.100 54.100 ;
        RECT 18.900 53.400 20.200 53.700 ;
        RECT 10.200 51.500 10.600 52.500 ;
        RECT 12.300 51.500 12.700 53.000 ;
        RECT 15.800 52.800 16.700 53.100 ;
        RECT 18.100 52.800 18.600 53.100 ;
        RECT 16.300 51.100 16.700 52.800 ;
        RECT 18.200 51.100 18.600 52.800 ;
        RECT 19.800 51.100 20.200 53.400 ;
        RECT 20.600 52.400 21.000 53.200 ;
        RECT 21.500 52.200 21.800 53.800 ;
        RECT 21.400 51.100 21.800 52.200 ;
        RECT 23.000 53.600 25.100 53.900 ;
        RECT 25.600 53.800 26.600 54.200 ;
        RECT 23.000 52.500 23.300 53.600 ;
        RECT 25.600 53.500 25.900 53.800 ;
        RECT 25.500 53.300 25.900 53.500 ;
        RECT 27.800 53.400 28.200 54.200 ;
        RECT 25.100 53.200 25.900 53.300 ;
        RECT 24.600 53.000 25.900 53.200 ;
        RECT 28.600 53.100 29.000 59.900 ;
        RECT 29.400 55.800 29.800 56.600 ;
        RECT 30.200 56.200 30.600 59.900 ;
        RECT 31.100 56.200 31.500 56.300 ;
        RECT 30.200 55.900 31.500 56.200 ;
        RECT 32.400 55.900 33.200 59.900 ;
        RECT 34.200 56.200 34.600 56.300 ;
        RECT 35.000 56.200 35.400 59.900 ;
        RECT 34.200 55.900 35.400 56.200 ;
        RECT 31.700 55.200 32.100 55.300 ;
        RECT 32.700 55.200 33.000 55.900 ;
        RECT 31.300 54.900 32.100 55.200 ;
        RECT 31.300 54.800 31.700 54.900 ;
        RECT 32.600 54.800 33.000 55.200 ;
        RECT 32.000 54.300 32.400 54.400 ;
        RECT 31.000 54.200 32.400 54.300 ;
        RECT 30.200 54.000 32.400 54.200 ;
        RECT 32.700 54.200 33.000 54.800 ;
        RECT 30.200 53.900 31.300 54.000 ;
        RECT 32.700 53.900 33.200 54.200 ;
        RECT 30.200 53.800 31.000 53.900 ;
        RECT 31.100 53.400 31.500 53.500 ;
        RECT 30.200 53.100 31.500 53.400 ;
        RECT 31.800 53.200 32.600 53.600 ;
        RECT 24.600 52.800 25.500 53.000 ;
        RECT 28.600 52.800 29.500 53.100 ;
        RECT 23.000 51.500 23.400 52.500 ;
        RECT 25.100 51.500 25.500 52.800 ;
        RECT 29.100 51.100 29.500 52.800 ;
        RECT 30.200 51.100 30.600 53.100 ;
        RECT 32.900 52.900 33.200 53.900 ;
        RECT 33.600 53.800 34.000 54.200 ;
        RECT 34.600 53.800 35.400 54.200 ;
        RECT 36.600 54.100 37.000 59.900 ;
        RECT 38.700 56.200 39.100 59.900 ;
        RECT 39.400 56.800 39.800 57.200 ;
        RECT 39.500 56.200 39.800 56.800 ;
        RECT 38.700 55.900 39.200 56.200 ;
        RECT 39.500 55.900 40.200 56.200 ;
        RECT 37.400 55.100 37.800 55.200 ;
        RECT 38.200 55.100 38.600 55.200 ;
        RECT 37.400 54.800 38.600 55.100 ;
        RECT 38.200 54.400 38.600 54.800 ;
        RECT 38.900 54.200 39.200 55.900 ;
        RECT 39.800 55.800 40.200 55.900 ;
        RECT 40.600 55.800 41.000 56.600 ;
        RECT 39.800 55.100 40.100 55.800 ;
        RECT 41.400 55.100 41.800 59.900 ;
        RECT 39.800 54.800 41.800 55.100 ;
        RECT 37.400 54.100 37.800 54.200 ;
        RECT 36.600 53.800 38.200 54.100 ;
        RECT 38.900 53.800 40.200 54.200 ;
        RECT 33.600 53.600 33.900 53.800 ;
        RECT 33.500 53.200 33.900 53.600 ;
        RECT 34.200 53.400 34.600 53.500 ;
        RECT 34.200 53.100 35.400 53.400 ;
        RECT 32.400 51.100 33.200 52.900 ;
        RECT 35.000 51.100 35.400 53.100 ;
        RECT 35.800 52.400 36.200 53.200 ;
        RECT 36.600 51.100 37.000 53.800 ;
        RECT 37.800 53.600 38.200 53.800 ;
        RECT 37.500 53.100 39.300 53.300 ;
        RECT 39.800 53.100 40.100 53.800 ;
        RECT 41.400 53.100 41.800 54.800 ;
        RECT 42.200 53.400 42.600 54.200 ;
        RECT 43.800 54.100 44.200 59.900 ;
        RECT 47.500 56.200 47.900 59.900 ;
        RECT 48.200 56.800 48.600 57.200 ;
        RECT 48.300 56.200 48.600 56.800 ;
        RECT 47.500 55.900 48.000 56.200 ;
        RECT 48.300 56.100 49.000 56.200 ;
        RECT 50.200 56.100 50.600 59.900 ;
        RECT 48.300 55.900 50.600 56.100 ;
        RECT 44.600 55.100 45.000 55.200 ;
        RECT 47.000 55.100 47.400 55.200 ;
        RECT 44.600 54.800 47.400 55.100 ;
        RECT 47.000 54.400 47.400 54.800 ;
        RECT 47.700 54.200 48.000 55.900 ;
        RECT 48.600 55.800 50.600 55.900 ;
        RECT 51.000 55.800 51.400 56.600 ;
        RECT 46.200 54.100 46.600 54.200 ;
        RECT 43.800 53.800 47.000 54.100 ;
        RECT 47.700 53.800 49.000 54.200 ;
        RECT 37.400 53.000 39.400 53.100 ;
        RECT 37.400 51.100 37.800 53.000 ;
        RECT 39.000 51.100 39.400 53.000 ;
        RECT 39.800 51.100 40.200 53.100 ;
        RECT 40.900 52.800 41.800 53.100 ;
        RECT 40.900 51.100 41.300 52.800 ;
        RECT 43.000 52.400 43.400 53.200 ;
        RECT 43.800 51.100 44.200 53.800 ;
        RECT 46.600 53.600 47.000 53.800 ;
        RECT 46.300 53.100 48.100 53.300 ;
        RECT 48.600 53.100 48.900 53.800 ;
        RECT 49.400 53.400 49.800 54.200 ;
        RECT 50.200 53.100 50.600 55.800 ;
        RECT 51.800 55.600 52.200 59.900 ;
        RECT 53.900 57.900 54.500 59.900 ;
        RECT 56.200 57.900 56.600 59.900 ;
        RECT 58.400 58.200 58.800 59.900 ;
        RECT 58.400 57.900 59.400 58.200 ;
        RECT 54.200 57.500 54.600 57.900 ;
        RECT 56.300 57.600 56.600 57.900 ;
        RECT 55.900 57.300 57.700 57.600 ;
        RECT 59.000 57.500 59.400 57.900 ;
        RECT 55.900 57.200 56.300 57.300 ;
        RECT 57.300 57.200 57.700 57.300 ;
        RECT 53.800 56.600 54.500 57.000 ;
        RECT 54.200 56.100 54.500 56.600 ;
        RECT 55.300 56.500 56.400 56.800 ;
        RECT 55.300 56.400 55.700 56.500 ;
        RECT 54.200 55.800 55.400 56.100 ;
        RECT 51.800 55.300 53.900 55.600 ;
        RECT 51.800 53.600 52.200 55.300 ;
        RECT 53.500 55.200 53.900 55.300 ;
        RECT 52.700 54.900 53.100 55.000 ;
        RECT 52.700 54.600 54.600 54.900 ;
        RECT 54.200 54.500 54.600 54.600 ;
        RECT 55.100 54.200 55.400 55.800 ;
        RECT 56.100 55.900 56.400 56.500 ;
        RECT 56.700 56.500 57.100 56.600 ;
        RECT 59.000 56.500 59.400 56.600 ;
        RECT 56.700 56.200 59.400 56.500 ;
        RECT 56.100 55.700 58.500 55.900 ;
        RECT 60.600 55.700 61.000 59.900 ;
        RECT 56.100 55.600 61.000 55.700 ;
        RECT 58.100 55.500 61.000 55.600 ;
        RECT 58.200 55.400 61.000 55.500 ;
        RECT 61.400 55.600 61.800 59.900 ;
        RECT 63.500 57.900 64.100 59.900 ;
        RECT 65.800 57.900 66.200 59.900 ;
        RECT 68.000 58.200 68.400 59.900 ;
        RECT 68.000 57.900 69.000 58.200 ;
        RECT 63.800 57.500 64.200 57.900 ;
        RECT 65.900 57.600 66.200 57.900 ;
        RECT 65.500 57.300 67.300 57.600 ;
        RECT 68.600 57.500 69.000 57.900 ;
        RECT 65.500 57.200 65.900 57.300 ;
        RECT 66.900 57.200 67.300 57.300 ;
        RECT 63.400 56.600 64.100 57.000 ;
        RECT 63.800 56.100 64.100 56.600 ;
        RECT 64.900 56.500 66.000 56.800 ;
        RECT 64.900 56.400 65.300 56.500 ;
        RECT 63.800 55.800 65.000 56.100 ;
        RECT 61.400 55.300 63.500 55.600 ;
        RECT 57.400 55.100 57.800 55.200 ;
        RECT 57.400 54.800 59.900 55.100 ;
        RECT 58.200 54.700 58.600 54.800 ;
        RECT 59.500 54.700 59.900 54.800 ;
        RECT 58.700 54.200 59.100 54.300 ;
        RECT 55.100 53.900 60.600 54.200 ;
        RECT 55.300 53.800 55.700 53.900 ;
        RECT 57.400 53.800 57.800 53.900 ;
        RECT 51.800 53.300 53.700 53.600 ;
        RECT 46.200 53.000 48.200 53.100 ;
        RECT 46.200 51.100 46.600 53.000 ;
        RECT 47.800 51.100 48.200 53.000 ;
        RECT 48.600 51.100 49.000 53.100 ;
        RECT 50.200 52.800 51.100 53.100 ;
        RECT 50.700 51.100 51.100 52.800 ;
        RECT 51.800 51.100 52.200 53.300 ;
        RECT 53.300 53.200 53.700 53.300 ;
        RECT 58.200 52.800 58.500 53.900 ;
        RECT 59.800 53.800 60.600 53.900 ;
        RECT 61.400 53.600 61.800 55.300 ;
        RECT 63.100 55.200 63.500 55.300 ;
        RECT 64.700 55.200 65.000 55.800 ;
        RECT 65.700 55.900 66.000 56.500 ;
        RECT 66.300 56.500 66.700 56.600 ;
        RECT 68.600 56.500 69.000 56.600 ;
        RECT 66.300 56.200 69.000 56.500 ;
        RECT 65.700 55.700 68.100 55.900 ;
        RECT 70.200 55.700 70.600 59.900 ;
        RECT 72.300 56.300 72.700 59.900 ;
        RECT 74.700 56.300 75.100 59.900 ;
        RECT 71.800 55.900 72.700 56.300 ;
        RECT 74.200 55.900 75.100 56.300 ;
        RECT 75.800 57.500 76.200 59.500 ;
        RECT 65.700 55.600 70.600 55.700 ;
        RECT 67.700 55.500 70.600 55.600 ;
        RECT 67.800 55.400 70.600 55.500 ;
        RECT 62.300 54.900 62.700 55.000 ;
        RECT 62.300 54.600 64.200 54.900 ;
        RECT 64.600 54.800 65.000 55.200 ;
        RECT 67.000 55.100 67.400 55.200 ;
        RECT 71.900 55.100 72.200 55.900 ;
        RECT 67.000 54.800 69.500 55.100 ;
        RECT 63.800 54.500 64.200 54.600 ;
        RECT 64.700 54.200 65.000 54.800 ;
        RECT 67.800 54.700 68.200 54.800 ;
        RECT 69.100 54.700 69.500 54.800 ;
        RECT 71.000 54.800 72.200 55.100 ;
        RECT 72.600 54.800 73.000 55.600 ;
        RECT 68.300 54.200 68.700 54.300 ;
        RECT 71.000 54.200 71.300 54.800 ;
        RECT 71.900 54.200 72.200 54.800 ;
        RECT 74.300 54.200 74.600 55.900 ;
        RECT 75.800 55.800 76.100 57.500 ;
        RECT 77.900 56.400 78.300 59.900 ;
        RECT 77.900 56.100 78.700 56.400 ;
        RECT 75.000 54.800 75.400 55.600 ;
        RECT 75.800 55.500 77.700 55.800 ;
        RECT 75.800 54.400 76.200 55.200 ;
        RECT 76.600 54.400 77.000 55.200 ;
        RECT 77.400 54.500 77.700 55.500 ;
        RECT 64.700 53.900 70.200 54.200 ;
        RECT 64.900 53.800 65.300 53.900 ;
        RECT 57.300 52.700 57.700 52.800 ;
        RECT 54.200 52.100 54.600 52.500 ;
        RECT 56.300 52.400 57.700 52.700 ;
        RECT 58.200 52.400 58.600 52.800 ;
        RECT 56.300 52.100 56.600 52.400 ;
        RECT 59.000 52.100 59.400 52.500 ;
        RECT 53.900 51.800 54.600 52.100 ;
        RECT 53.900 51.100 54.500 51.800 ;
        RECT 56.200 51.100 56.600 52.100 ;
        RECT 58.400 51.800 59.400 52.100 ;
        RECT 58.400 51.100 58.800 51.800 ;
        RECT 60.600 51.100 61.000 53.500 ;
        RECT 61.400 53.300 63.300 53.600 ;
        RECT 61.400 51.100 61.800 53.300 ;
        RECT 62.900 53.200 63.300 53.300 ;
        RECT 67.800 52.800 68.100 53.900 ;
        RECT 69.400 53.800 70.200 53.900 ;
        RECT 71.000 53.800 71.400 54.200 ;
        RECT 71.800 53.800 72.200 54.200 ;
        RECT 74.200 53.800 74.600 54.200 ;
        RECT 77.400 54.100 78.100 54.500 ;
        RECT 78.400 54.200 78.700 56.100 ;
        RECT 80.600 56.200 81.000 59.900 ;
        RECT 82.200 59.600 84.200 59.900 ;
        RECT 82.200 56.200 82.600 59.600 ;
        RECT 80.600 55.900 82.600 56.200 ;
        RECT 83.000 55.800 83.400 59.300 ;
        RECT 83.800 55.900 84.200 59.600 ;
        RECT 84.600 55.900 85.000 59.900 ;
        RECT 85.400 56.200 85.800 59.900 ;
        RECT 87.000 56.200 87.400 59.900 ;
        RECT 89.100 56.300 89.500 59.900 ;
        RECT 85.400 55.900 87.400 56.200 ;
        RECT 88.600 55.900 89.500 56.300 ;
        RECT 83.000 55.600 83.300 55.800 ;
        RECT 79.000 54.800 79.400 55.600 ;
        RECT 81.000 55.200 81.400 55.400 ;
        RECT 82.300 55.300 83.300 55.600 ;
        RECT 82.300 55.200 82.600 55.300 ;
        RECT 80.600 54.900 81.400 55.200 ;
        RECT 80.600 54.800 81.000 54.900 ;
        RECT 82.200 54.800 82.600 55.200 ;
        RECT 83.800 54.800 84.200 55.600 ;
        RECT 84.700 55.200 85.000 55.900 ;
        RECT 86.600 55.200 87.000 55.400 ;
        RECT 88.700 55.200 89.000 55.900 ;
        RECT 84.600 54.900 85.800 55.200 ;
        RECT 86.600 54.900 87.400 55.200 ;
        RECT 84.600 54.800 85.000 54.900 ;
        RECT 77.400 53.900 77.900 54.100 ;
        RECT 66.900 52.700 67.300 52.800 ;
        RECT 63.800 52.100 64.200 52.500 ;
        RECT 65.900 52.400 67.300 52.700 ;
        RECT 67.800 52.400 68.200 52.800 ;
        RECT 65.900 52.100 66.200 52.400 ;
        RECT 68.600 52.100 69.000 52.500 ;
        RECT 63.500 51.800 64.200 52.100 ;
        RECT 63.500 51.100 64.100 51.800 ;
        RECT 65.800 51.100 66.200 52.100 ;
        RECT 68.000 51.800 69.000 52.100 ;
        RECT 68.000 51.100 68.400 51.800 ;
        RECT 70.200 51.100 70.600 53.500 ;
        RECT 71.000 52.400 71.400 53.200 ;
        RECT 71.900 52.100 72.200 53.800 ;
        RECT 73.400 52.400 73.800 53.200 ;
        RECT 74.300 52.200 74.600 53.800 ;
        RECT 71.800 51.100 72.200 52.100 ;
        RECT 74.200 51.100 74.600 52.200 ;
        RECT 75.800 53.600 77.900 53.900 ;
        RECT 78.400 53.800 79.400 54.200 ;
        RECT 81.400 53.800 81.800 54.600 ;
        RECT 75.800 52.500 76.100 53.600 ;
        RECT 78.400 53.500 78.700 53.800 ;
        RECT 78.300 53.300 78.700 53.500 ;
        RECT 77.900 53.200 78.700 53.300 ;
        RECT 77.400 53.000 78.700 53.200 ;
        RECT 82.300 53.100 82.600 54.800 ;
        RECT 82.900 54.400 83.300 54.800 ;
        RECT 83.000 54.200 83.300 54.400 ;
        RECT 83.000 53.800 83.400 54.200 ;
        RECT 77.400 52.800 78.300 53.000 ;
        RECT 75.800 51.500 76.200 52.500 ;
        RECT 77.900 51.500 78.300 52.800 ;
        RECT 82.100 51.100 82.900 53.100 ;
        RECT 84.600 52.800 85.000 53.200 ;
        RECT 85.500 53.100 85.800 54.900 ;
        RECT 87.000 54.800 87.400 54.900 ;
        RECT 88.600 54.800 89.000 55.200 ;
        RECT 89.400 55.100 89.800 55.600 ;
        RECT 91.000 55.100 91.400 59.900 ;
        RECT 91.800 56.100 92.200 56.600 ;
        RECT 93.400 56.100 93.800 59.900 ;
        RECT 95.800 56.900 96.200 59.900 ;
        RECT 95.900 56.600 96.200 56.900 ;
        RECT 97.400 59.600 99.400 59.900 ;
        RECT 97.400 56.900 97.800 59.600 ;
        RECT 98.200 56.900 98.600 59.300 ;
        RECT 99.000 57.000 99.400 59.600 ;
        RECT 99.900 59.600 101.700 59.900 ;
        RECT 99.900 59.500 100.200 59.600 ;
        RECT 97.400 56.600 97.700 56.900 ;
        RECT 95.900 56.300 97.700 56.600 ;
        RECT 98.300 56.700 98.600 56.900 ;
        RECT 99.800 56.700 100.200 59.500 ;
        RECT 101.400 59.500 101.700 59.600 ;
        RECT 98.300 56.500 100.200 56.700 ;
        RECT 100.600 56.500 101.000 59.300 ;
        RECT 101.400 56.500 101.800 59.500 ;
        RECT 98.300 56.400 100.100 56.500 ;
        RECT 100.600 56.200 100.900 56.500 ;
        RECT 102.200 56.200 102.600 59.900 ;
        RECT 103.800 59.600 105.800 59.900 ;
        RECT 103.800 56.200 104.200 59.600 ;
        RECT 100.600 56.100 101.000 56.200 ;
        RECT 91.800 55.800 93.800 56.100 ;
        RECT 89.400 54.800 91.400 55.100 ;
        RECT 86.200 53.800 86.600 54.600 ;
        RECT 88.700 54.200 89.000 54.800 ;
        RECT 88.600 53.800 89.000 54.200 ;
        RECT 84.700 52.400 85.100 52.800 ;
        RECT 85.400 51.100 85.800 53.100 ;
        RECT 87.800 52.400 88.200 53.200 ;
        RECT 88.700 52.100 89.000 53.800 ;
        RECT 90.200 53.400 90.600 54.200 ;
        RECT 91.000 53.100 91.400 54.800 ;
        RECT 93.400 55.100 93.800 55.800 ;
        RECT 99.300 55.800 101.000 56.100 ;
        RECT 102.200 55.900 104.200 56.200 ;
        RECT 104.600 55.900 105.000 59.300 ;
        RECT 105.400 55.900 105.800 59.600 ;
        RECT 106.500 56.300 106.900 59.900 ;
        RECT 109.400 57.900 109.800 59.900 ;
        RECT 106.500 55.900 107.400 56.300 ;
        RECT 98.200 55.100 99.000 55.200 ;
        RECT 93.400 54.800 99.000 55.100 ;
        RECT 91.000 52.800 91.900 53.100 ;
        RECT 88.600 51.100 89.000 52.100 ;
        RECT 91.500 51.100 91.900 52.800 ;
        RECT 92.600 52.400 93.000 53.200 ;
        RECT 93.400 51.100 93.800 54.800 ;
        RECT 95.800 54.100 96.200 54.200 ;
        RECT 97.400 54.100 98.200 54.200 ;
        RECT 95.800 53.800 98.200 54.100 ;
        RECT 95.000 53.100 95.400 53.200 ;
        RECT 96.600 53.100 97.500 53.200 ;
        RECT 95.000 52.800 97.500 53.100 ;
        RECT 99.300 52.500 99.600 55.800 ;
        RECT 104.600 55.600 104.900 55.900 ;
        RECT 102.600 55.200 103.000 55.400 ;
        RECT 103.900 55.300 104.900 55.600 ;
        RECT 103.900 55.200 104.200 55.300 ;
        RECT 102.200 54.900 103.000 55.200 ;
        RECT 102.200 54.800 102.600 54.900 ;
        RECT 103.800 54.800 104.200 55.200 ;
        RECT 105.400 54.800 105.800 55.600 ;
        RECT 106.200 54.800 106.600 55.600 ;
        RECT 103.000 53.800 103.400 54.600 ;
        RECT 103.900 53.100 104.200 54.800 ;
        RECT 104.500 54.400 104.900 54.800 ;
        RECT 104.600 54.200 104.900 54.400 ;
        RECT 107.000 54.200 107.300 55.900 ;
        RECT 109.500 55.800 109.800 57.900 ;
        RECT 111.000 55.900 111.400 59.900 ;
        RECT 111.800 59.600 113.800 59.900 ;
        RECT 111.800 55.900 112.200 59.600 ;
        RECT 112.600 55.900 113.000 59.300 ;
        RECT 113.400 56.200 113.800 59.600 ;
        RECT 115.000 56.200 115.400 59.900 ;
        RECT 116.100 56.200 116.500 59.900 ;
        RECT 113.400 55.900 115.400 56.200 ;
        RECT 115.800 55.900 116.500 56.200 ;
        RECT 109.500 55.500 110.700 55.800 ;
        RECT 107.800 55.100 108.200 55.200 ;
        RECT 107.800 54.800 109.000 55.100 ;
        RECT 109.400 54.800 109.800 55.200 ;
        RECT 104.600 54.100 105.000 54.200 ;
        RECT 107.000 54.100 107.400 54.200 ;
        RECT 108.600 54.100 109.000 54.800 ;
        RECT 109.500 54.400 109.800 54.800 ;
        RECT 109.500 54.100 110.000 54.400 ;
        RECT 104.600 53.800 109.000 54.100 ;
        RECT 109.600 54.000 110.000 54.100 ;
        RECT 110.400 53.800 110.700 55.500 ;
        RECT 111.100 55.200 111.400 55.900 ;
        RECT 112.700 55.600 113.000 55.900 ;
        RECT 115.800 55.800 116.200 55.900 ;
        RECT 111.000 54.800 111.400 55.200 ;
        RECT 111.800 54.800 112.200 55.600 ;
        RECT 112.700 55.300 113.700 55.600 ;
        RECT 113.400 55.200 113.700 55.300 ;
        RECT 114.600 55.200 115.000 55.400 ;
        RECT 115.800 55.200 116.100 55.800 ;
        RECT 118.200 55.600 118.600 59.900 ;
        RECT 119.000 56.200 119.400 59.900 ;
        RECT 120.600 56.200 121.000 59.900 ;
        RECT 119.000 55.900 121.000 56.200 ;
        RECT 121.400 55.900 121.800 59.900 ;
        RECT 122.200 56.200 122.600 59.900 ;
        RECT 122.200 55.900 123.300 56.200 ;
        RECT 123.800 55.900 124.200 59.900 ;
        RECT 116.600 55.400 118.600 55.600 ;
        RECT 116.500 55.300 118.600 55.400 ;
        RECT 113.400 54.800 113.800 55.200 ;
        RECT 114.600 54.900 115.400 55.200 ;
        RECT 115.000 54.800 115.400 54.900 ;
        RECT 115.800 54.800 116.200 55.200 ;
        RECT 116.500 55.000 116.900 55.300 ;
        RECT 119.400 55.200 119.800 55.400 ;
        RECT 121.400 55.200 121.700 55.900 ;
        RECT 123.000 55.600 123.300 55.900 ;
        RECT 123.000 55.200 123.600 55.600 ;
        RECT 97.600 52.200 99.600 52.500 ;
        RECT 97.400 51.800 97.900 52.200 ;
        RECT 99.000 52.100 99.600 52.200 ;
        RECT 101.400 52.100 101.800 52.200 ;
        RECT 99.000 51.800 101.800 52.100 ;
        RECT 97.400 51.100 97.800 51.800 ;
        RECT 99.000 51.100 99.400 51.800 ;
        RECT 103.700 51.100 104.500 53.100 ;
        RECT 107.000 52.100 107.300 53.800 ;
        RECT 110.400 53.700 110.800 53.800 ;
        RECT 109.300 53.500 110.800 53.700 ;
        RECT 108.700 53.400 110.800 53.500 ;
        RECT 108.700 53.200 109.600 53.400 ;
        RECT 107.800 52.400 108.200 53.200 ;
        RECT 108.700 53.100 109.000 53.200 ;
        RECT 111.100 53.100 111.400 54.800 ;
        RECT 112.700 54.400 113.100 54.800 ;
        RECT 112.700 54.200 113.000 54.400 ;
        RECT 112.600 53.800 113.000 54.200 ;
        RECT 113.400 53.100 113.700 54.800 ;
        RECT 114.200 53.800 114.600 54.600 ;
        RECT 115.800 53.100 116.100 54.800 ;
        RECT 116.500 53.500 116.800 55.000 ;
        RECT 119.000 54.900 119.800 55.200 ;
        RECT 120.600 54.900 121.800 55.200 ;
        RECT 119.000 54.800 119.400 54.900 ;
        RECT 117.200 54.200 117.600 54.600 ;
        RECT 117.300 53.800 117.800 54.200 ;
        RECT 119.000 54.100 119.400 54.200 ;
        RECT 119.800 54.100 120.200 54.600 ;
        RECT 119.000 53.800 120.200 54.100 ;
        RECT 120.600 54.100 120.900 54.900 ;
        RECT 121.400 54.800 121.800 54.900 ;
        RECT 122.200 54.400 122.600 55.200 ;
        RECT 121.400 54.100 121.800 54.200 ;
        RECT 120.600 53.800 121.800 54.100 ;
        RECT 116.500 53.200 117.700 53.500 ;
        RECT 107.000 51.100 107.400 52.100 ;
        RECT 108.600 51.100 109.000 53.100 ;
        RECT 110.700 52.600 111.400 53.100 ;
        RECT 110.700 51.100 111.100 52.600 ;
        RECT 113.100 51.100 113.900 53.100 ;
        RECT 115.800 51.100 116.200 53.100 ;
        RECT 117.400 52.100 117.700 53.200 ;
        RECT 118.200 52.400 118.600 53.200 ;
        RECT 120.600 53.100 120.900 53.800 ;
        RECT 123.000 53.700 123.300 55.200 ;
        RECT 123.900 54.800 124.200 55.900 ;
        RECT 122.200 53.400 123.300 53.700 ;
        RECT 117.400 51.100 117.800 52.100 ;
        RECT 120.600 51.100 121.000 53.100 ;
        RECT 121.400 52.800 121.800 53.200 ;
        RECT 121.300 52.400 121.700 52.800 ;
        RECT 122.200 51.100 122.600 53.400 ;
        RECT 123.800 51.100 124.200 54.800 ;
        RECT 124.600 55.600 125.000 59.900 ;
        RECT 126.700 57.900 127.300 59.900 ;
        RECT 129.000 57.900 129.400 59.900 ;
        RECT 131.200 58.200 131.600 59.900 ;
        RECT 131.200 57.900 132.200 58.200 ;
        RECT 127.000 57.500 127.400 57.900 ;
        RECT 129.100 57.600 129.400 57.900 ;
        RECT 128.700 57.300 130.500 57.600 ;
        RECT 131.800 57.500 132.200 57.900 ;
        RECT 128.700 57.200 129.100 57.300 ;
        RECT 130.100 57.200 130.500 57.300 ;
        RECT 126.600 56.600 127.300 57.000 ;
        RECT 127.000 56.100 127.300 56.600 ;
        RECT 128.100 56.500 129.200 56.800 ;
        RECT 128.100 56.400 128.500 56.500 ;
        RECT 127.000 55.800 128.200 56.100 ;
        RECT 124.600 55.300 126.700 55.600 ;
        RECT 124.600 53.600 125.000 55.300 ;
        RECT 126.300 55.200 126.700 55.300 ;
        RECT 125.500 54.900 125.900 55.000 ;
        RECT 125.500 54.600 127.400 54.900 ;
        RECT 127.000 54.500 127.400 54.600 ;
        RECT 127.900 54.200 128.200 55.800 ;
        RECT 128.900 55.900 129.200 56.500 ;
        RECT 129.500 56.500 129.900 56.600 ;
        RECT 131.800 56.500 132.200 56.600 ;
        RECT 129.500 56.200 132.200 56.500 ;
        RECT 128.900 55.700 131.300 55.900 ;
        RECT 133.400 55.700 133.800 59.900 ;
        RECT 134.200 55.900 134.600 59.900 ;
        RECT 135.000 56.200 135.400 59.900 ;
        RECT 136.600 56.200 137.000 59.900 ;
        RECT 135.000 55.900 137.000 56.200 ;
        RECT 137.400 55.900 137.800 59.900 ;
        RECT 138.200 56.200 138.600 59.900 ;
        RECT 139.800 56.200 140.200 59.900 ;
        RECT 138.200 55.900 140.200 56.200 ;
        RECT 128.900 55.600 133.800 55.700 ;
        RECT 130.900 55.500 133.800 55.600 ;
        RECT 131.000 55.400 133.800 55.500 ;
        RECT 134.300 55.200 134.600 55.900 ;
        RECT 136.200 55.200 136.600 55.400 ;
        RECT 137.500 55.200 137.800 55.900 ;
        RECT 139.400 55.200 139.800 55.400 ;
        RECT 130.200 55.100 130.600 55.200 ;
        RECT 130.200 54.800 132.700 55.100 ;
        RECT 134.200 54.900 135.400 55.200 ;
        RECT 136.200 54.900 137.000 55.200 ;
        RECT 134.200 54.800 134.600 54.900 ;
        RECT 132.300 54.700 132.700 54.800 ;
        RECT 131.500 54.200 131.900 54.300 ;
        RECT 127.800 54.100 133.400 54.200 ;
        RECT 127.800 53.900 134.500 54.100 ;
        RECT 127.800 53.800 128.500 53.900 ;
        RECT 129.400 53.800 129.800 53.900 ;
        RECT 124.600 53.300 126.500 53.600 ;
        RECT 124.600 51.100 125.000 53.300 ;
        RECT 126.100 53.200 126.500 53.300 ;
        RECT 131.000 52.800 131.300 53.900 ;
        RECT 132.600 53.800 134.500 53.900 ;
        RECT 130.100 52.700 130.500 52.800 ;
        RECT 127.000 52.100 127.400 52.500 ;
        RECT 129.100 52.400 130.500 52.700 ;
        RECT 131.000 52.400 131.400 52.800 ;
        RECT 129.100 52.100 129.400 52.400 ;
        RECT 131.800 52.100 132.200 52.500 ;
        RECT 126.700 51.800 127.400 52.100 ;
        RECT 126.700 51.100 127.300 51.800 ;
        RECT 129.000 51.100 129.400 52.100 ;
        RECT 131.200 51.800 132.200 52.100 ;
        RECT 131.200 51.100 131.600 51.800 ;
        RECT 133.400 51.100 133.800 53.500 ;
        RECT 134.200 53.200 134.500 53.800 ;
        RECT 134.200 52.800 134.600 53.200 ;
        RECT 135.100 53.100 135.400 54.900 ;
        RECT 136.600 54.800 137.000 54.900 ;
        RECT 137.400 54.900 138.600 55.200 ;
        RECT 139.400 54.900 140.200 55.200 ;
        RECT 137.400 54.800 137.800 54.900 ;
        RECT 135.800 54.100 136.200 54.600 ;
        RECT 138.300 54.100 138.600 54.900 ;
        RECT 139.800 54.800 140.200 54.900 ;
        RECT 135.800 53.800 138.600 54.100 ;
        RECT 139.000 53.800 139.400 54.600 ;
        RECT 141.400 54.100 141.800 59.900 ;
        RECT 142.200 54.100 142.600 54.200 ;
        RECT 141.400 53.800 142.600 54.100 ;
        RECT 134.300 52.400 134.700 52.800 ;
        RECT 135.000 51.100 135.400 53.100 ;
        RECT 137.400 52.800 137.800 53.200 ;
        RECT 138.300 53.100 138.600 53.800 ;
        RECT 137.500 52.400 137.900 52.800 ;
        RECT 138.200 51.100 138.600 53.100 ;
        RECT 140.600 52.400 141.000 53.200 ;
        RECT 141.400 51.100 141.800 53.800 ;
        RECT 142.200 53.400 142.600 53.800 ;
        RECT 143.000 54.100 143.400 59.900 ;
        RECT 143.800 55.800 144.200 56.600 ;
        RECT 144.600 56.200 145.000 59.900 ;
        RECT 146.200 56.200 146.600 59.900 ;
        RECT 144.600 55.900 146.600 56.200 ;
        RECT 147.000 55.900 147.400 59.900 ;
        RECT 149.800 56.800 150.200 57.200 ;
        RECT 149.800 56.200 150.100 56.800 ;
        RECT 150.500 56.200 150.900 59.900 ;
        RECT 149.400 55.900 150.100 56.200 ;
        RECT 150.400 55.900 150.900 56.200 ;
        RECT 145.000 55.200 145.400 55.400 ;
        RECT 147.000 55.200 147.300 55.900 ;
        RECT 149.400 55.800 149.800 55.900 ;
        RECT 144.600 54.900 145.400 55.200 ;
        RECT 146.200 54.900 147.400 55.200 ;
        RECT 144.600 54.800 145.000 54.900 ;
        RECT 145.400 54.100 145.800 54.600 ;
        RECT 143.000 53.800 145.800 54.100 ;
        RECT 143.000 53.100 143.400 53.800 ;
        RECT 146.200 53.100 146.500 54.900 ;
        RECT 147.000 54.800 147.400 54.900 ;
        RECT 150.400 54.200 150.700 55.900 ;
        RECT 151.000 55.100 151.400 55.200 ;
        RECT 153.400 55.100 153.800 59.900 ;
        RECT 154.200 56.200 154.600 59.900 ;
        RECT 155.000 56.200 155.400 56.300 ;
        RECT 156.400 56.200 157.200 59.900 ;
        RECT 154.200 55.900 155.400 56.200 ;
        RECT 156.200 55.900 157.200 56.200 ;
        RECT 158.300 56.200 158.700 56.300 ;
        RECT 159.000 56.200 159.400 59.900 ;
        RECT 158.300 55.900 159.400 56.200 ;
        RECT 160.100 56.300 160.500 59.900 ;
        RECT 162.200 57.900 162.600 59.900 ;
        RECT 162.300 57.800 162.600 57.900 ;
        RECT 163.800 57.900 164.200 59.900 ;
        RECT 163.800 57.800 164.100 57.900 ;
        RECT 162.300 57.500 164.100 57.800 ;
        RECT 160.100 55.900 161.000 56.300 ;
        RECT 162.300 56.200 162.600 57.500 ;
        RECT 163.000 56.400 163.400 57.200 ;
        RECT 156.200 55.200 156.500 55.900 ;
        RECT 158.300 55.600 158.600 55.900 ;
        RECT 160.600 55.800 161.000 55.900 ;
        RECT 162.200 55.800 162.600 56.200 ;
        RECT 156.900 55.300 158.600 55.600 ;
        RECT 156.900 55.200 157.300 55.300 ;
        RECT 151.000 54.800 153.800 55.100 ;
        RECT 155.800 54.900 156.500 55.200 ;
        RECT 159.000 55.100 159.400 55.200 ;
        RECT 159.800 55.100 160.200 55.600 ;
        RECT 158.000 54.900 158.400 55.000 ;
        RECT 155.800 54.800 156.700 54.900 ;
        RECT 151.000 54.400 151.400 54.800 ;
        RECT 147.000 54.100 147.400 54.200 ;
        RECT 149.400 54.100 150.700 54.200 ;
        RECT 151.800 54.100 152.200 54.200 ;
        RECT 147.000 53.800 150.700 54.100 ;
        RECT 151.400 53.800 152.200 54.100 ;
        RECT 147.000 53.100 147.400 53.200 ;
        RECT 147.800 53.100 148.200 53.200 ;
        RECT 149.500 53.100 149.800 53.800 ;
        RECT 151.400 53.600 151.800 53.800 ;
        RECT 152.600 53.400 153.000 54.200 ;
        RECT 153.400 54.100 153.800 54.800 ;
        RECT 156.200 54.600 156.700 54.800 ;
        RECT 154.200 54.100 155.000 54.200 ;
        RECT 153.400 53.800 155.000 54.100 ;
        RECT 155.600 53.800 156.000 54.200 ;
        RECT 150.300 53.100 152.100 53.300 ;
        RECT 143.000 52.800 143.900 53.100 ;
        RECT 143.500 51.100 143.900 52.800 ;
        RECT 146.200 51.100 146.600 53.100 ;
        RECT 147.000 52.800 148.200 53.100 ;
        RECT 146.900 52.400 147.300 52.800 ;
        RECT 149.400 51.100 149.800 53.100 ;
        RECT 150.200 53.000 152.200 53.100 ;
        RECT 150.200 51.100 150.600 53.000 ;
        RECT 151.800 51.100 152.200 53.000 ;
        RECT 153.400 51.100 153.800 53.800 ;
        RECT 155.700 53.600 156.000 53.800 ;
        RECT 155.000 53.400 155.400 53.500 ;
        RECT 154.200 53.100 155.400 53.400 ;
        RECT 155.700 53.200 156.100 53.600 ;
        RECT 154.200 51.100 154.600 53.100 ;
        RECT 156.400 52.900 156.700 54.600 ;
        RECT 157.100 54.600 158.400 54.900 ;
        RECT 159.000 54.800 160.200 55.100 ;
        RECT 157.100 54.300 157.400 54.600 ;
        RECT 157.000 53.900 157.400 54.300 ;
        RECT 160.600 54.200 160.900 55.800 ;
        RECT 162.300 54.200 162.600 55.800 ;
        RECT 163.400 54.800 164.200 55.200 ;
        RECT 164.600 54.800 165.000 56.200 ;
        RECT 158.600 54.100 159.400 54.200 ;
        RECT 157.700 53.800 159.400 54.100 ;
        RECT 160.600 53.800 161.000 54.200 ;
        RECT 161.400 53.800 161.800 54.200 ;
        RECT 162.300 54.100 163.100 54.200 ;
        RECT 162.300 53.900 163.200 54.100 ;
        RECT 157.700 53.600 158.000 53.800 ;
        RECT 157.000 53.300 158.000 53.600 ;
        RECT 158.300 53.400 158.700 53.500 ;
        RECT 157.000 53.200 157.800 53.300 ;
        RECT 158.300 53.100 159.400 53.400 ;
        RECT 156.400 52.200 157.200 52.900 ;
        RECT 155.800 51.800 157.200 52.200 ;
        RECT 156.400 51.100 157.200 51.800 ;
        RECT 159.000 51.100 159.400 53.100 ;
        RECT 160.600 52.100 160.900 53.800 ;
        RECT 161.400 53.200 161.700 53.800 ;
        RECT 161.400 52.400 161.800 53.200 ;
        RECT 160.600 51.100 161.000 52.100 ;
        RECT 162.800 51.100 163.200 53.900 ;
        RECT 165.400 53.400 165.800 54.200 ;
        RECT 166.200 53.100 166.600 59.900 ;
        RECT 167.000 55.800 167.400 56.600 ;
        RECT 169.100 56.300 169.500 59.900 ;
        RECT 171.000 57.800 171.400 59.900 ;
        RECT 172.600 57.900 173.000 59.900 ;
        RECT 172.600 57.800 172.900 57.900 ;
        RECT 171.100 57.500 172.900 57.800 ;
        RECT 171.800 56.400 172.200 57.200 ;
        RECT 168.600 55.900 169.500 56.300 ;
        RECT 172.600 56.200 172.900 57.500 ;
        RECT 168.700 54.200 169.000 55.900 ;
        RECT 169.400 54.800 169.800 55.600 ;
        RECT 170.200 55.400 170.600 56.200 ;
        RECT 172.600 55.800 173.000 56.200 ;
        RECT 174.200 56.100 174.600 59.900 ;
        RECT 175.400 56.800 175.800 57.200 ;
        RECT 175.400 56.200 175.700 56.800 ;
        RECT 176.100 56.200 176.500 59.900 ;
        RECT 179.500 56.300 179.900 59.900 ;
        RECT 175.000 56.100 175.700 56.200 ;
        RECT 174.200 55.900 175.700 56.100 ;
        RECT 176.000 55.900 176.500 56.200 ;
        RECT 179.000 55.900 179.900 56.300 ;
        RECT 181.000 56.800 181.400 57.200 ;
        RECT 181.000 56.200 181.300 56.800 ;
        RECT 181.700 56.200 182.100 59.900 ;
        RECT 180.600 55.900 181.300 56.200 ;
        RECT 181.600 55.900 182.100 56.200 ;
        RECT 174.200 55.800 175.400 55.900 ;
        RECT 171.000 54.800 171.800 55.200 ;
        RECT 172.600 54.200 172.900 55.800 ;
        RECT 168.600 53.800 169.000 54.200 ;
        RECT 172.100 54.100 172.900 54.200 ;
        RECT 167.800 53.100 168.200 53.200 ;
        RECT 166.200 52.800 168.200 53.100 ;
        RECT 166.700 51.100 167.100 52.800 ;
        RECT 167.800 52.400 168.200 52.800 ;
        RECT 168.700 52.200 169.000 53.800 ;
        RECT 168.600 51.100 169.000 52.200 ;
        RECT 172.000 53.900 172.900 54.100 ;
        RECT 172.000 51.100 172.400 53.900 ;
        RECT 173.400 52.400 173.800 53.200 ;
        RECT 174.200 51.100 174.600 55.800 ;
        RECT 175.000 55.100 175.400 55.200 ;
        RECT 176.000 55.100 176.300 55.900 ;
        RECT 175.000 54.800 176.300 55.100 ;
        RECT 176.000 54.200 176.300 54.800 ;
        RECT 176.600 54.400 177.000 55.200 ;
        RECT 179.100 54.200 179.400 55.900 ;
        RECT 180.600 55.800 181.000 55.900 ;
        RECT 179.800 54.800 180.200 55.600 ;
        RECT 181.600 54.200 181.900 55.900 ;
        RECT 183.800 55.700 184.200 59.900 ;
        RECT 186.000 58.200 186.400 59.900 ;
        RECT 185.400 57.900 186.400 58.200 ;
        RECT 188.200 57.900 188.600 59.900 ;
        RECT 190.300 57.900 190.900 59.900 ;
        RECT 185.400 57.500 185.800 57.900 ;
        RECT 188.200 57.600 188.500 57.900 ;
        RECT 187.100 57.300 188.900 57.600 ;
        RECT 190.200 57.500 190.600 57.900 ;
        RECT 187.100 57.200 187.500 57.300 ;
        RECT 188.500 57.200 188.900 57.300 ;
        RECT 185.400 56.500 185.800 56.600 ;
        RECT 187.700 56.500 188.100 56.600 ;
        RECT 185.400 56.200 188.100 56.500 ;
        RECT 188.400 56.500 189.500 56.800 ;
        RECT 188.400 55.900 188.700 56.500 ;
        RECT 189.100 56.400 189.500 56.500 ;
        RECT 190.300 56.600 191.000 57.000 ;
        RECT 190.300 56.100 190.600 56.600 ;
        RECT 186.300 55.700 188.700 55.900 ;
        RECT 183.800 55.600 188.700 55.700 ;
        RECT 189.400 55.800 190.600 56.100 ;
        RECT 183.800 55.500 186.700 55.600 ;
        RECT 183.800 55.400 186.600 55.500 ;
        RECT 182.200 54.400 182.600 55.200 ;
        RECT 187.000 55.100 187.400 55.200 ;
        RECT 184.900 54.800 187.400 55.100 ;
        RECT 184.900 54.700 185.300 54.800 ;
        RECT 186.200 54.700 186.600 54.800 ;
        RECT 185.700 54.200 186.100 54.300 ;
        RECT 189.400 54.200 189.700 55.800 ;
        RECT 192.600 55.600 193.000 59.900 ;
        RECT 190.900 55.300 193.000 55.600 ;
        RECT 190.900 55.200 191.300 55.300 ;
        RECT 191.700 54.900 192.100 55.000 ;
        RECT 190.200 54.600 192.100 54.900 ;
        RECT 190.200 54.500 190.600 54.600 ;
        RECT 175.000 53.800 176.300 54.200 ;
        RECT 177.400 54.100 177.800 54.200 ;
        RECT 177.000 53.800 177.800 54.100 ;
        RECT 178.200 54.100 178.600 54.200 ;
        RECT 179.000 54.100 179.400 54.200 ;
        RECT 178.200 53.800 179.400 54.100 ;
        RECT 180.600 53.800 181.900 54.200 ;
        RECT 183.000 54.100 183.400 54.200 ;
        RECT 182.600 53.800 183.400 54.100 ;
        RECT 184.200 53.900 189.700 54.200 ;
        RECT 184.200 53.800 185.000 53.900 ;
        RECT 175.100 53.100 175.400 53.800 ;
        RECT 177.000 53.600 177.400 53.800 ;
        RECT 175.900 53.100 177.700 53.300 ;
        RECT 175.000 51.100 175.400 53.100 ;
        RECT 175.800 53.000 177.800 53.100 ;
        RECT 175.800 51.100 176.200 53.000 ;
        RECT 177.400 51.100 177.800 53.000 ;
        RECT 178.200 52.400 178.600 53.200 ;
        RECT 179.100 52.100 179.400 53.800 ;
        RECT 180.700 53.100 181.000 53.800 ;
        RECT 182.600 53.600 183.000 53.800 ;
        RECT 181.500 53.100 183.300 53.300 ;
        RECT 179.000 51.100 179.400 52.100 ;
        RECT 180.600 51.100 181.000 53.100 ;
        RECT 181.400 53.000 183.400 53.100 ;
        RECT 181.400 51.100 181.800 53.000 ;
        RECT 183.000 51.100 183.400 53.000 ;
        RECT 183.800 51.100 184.200 53.500 ;
        RECT 186.300 52.800 186.600 53.900 ;
        RECT 187.000 53.800 187.400 53.900 ;
        RECT 189.100 53.800 189.500 53.900 ;
        RECT 192.600 53.600 193.000 55.300 ;
        RECT 191.000 53.300 193.000 53.600 ;
        RECT 191.000 53.200 191.500 53.300 ;
        RECT 191.000 52.800 191.400 53.200 ;
        RECT 185.400 52.100 185.800 52.500 ;
        RECT 186.200 52.400 186.600 52.800 ;
        RECT 187.100 52.700 187.500 52.800 ;
        RECT 187.100 52.400 188.500 52.700 ;
        RECT 188.200 52.100 188.500 52.400 ;
        RECT 190.200 52.100 190.600 52.500 ;
        RECT 185.400 51.800 186.400 52.100 ;
        RECT 186.000 51.100 186.400 51.800 ;
        RECT 188.200 51.100 188.600 52.100 ;
        RECT 190.200 51.800 190.900 52.100 ;
        RECT 190.300 51.100 190.900 51.800 ;
        RECT 192.600 51.100 193.000 53.300 ;
        RECT 193.400 51.100 193.800 59.900 ;
        RECT 194.200 52.400 194.600 53.200 ;
        RECT 2.200 47.600 2.600 49.900 ;
        RECT 1.500 47.300 2.600 47.600 ;
        RECT 3.000 47.700 3.400 49.900 ;
        RECT 5.100 49.200 5.700 49.900 ;
        RECT 5.100 48.900 5.800 49.200 ;
        RECT 7.400 48.900 7.800 49.900 ;
        RECT 9.600 49.200 10.000 49.900 ;
        RECT 9.600 48.900 10.600 49.200 ;
        RECT 5.400 48.500 5.800 48.900 ;
        RECT 7.500 48.600 7.800 48.900 ;
        RECT 7.500 48.300 8.900 48.600 ;
        RECT 8.500 48.200 8.900 48.300 ;
        RECT 9.400 48.200 9.800 48.600 ;
        RECT 10.200 48.500 10.600 48.900 ;
        RECT 4.500 47.700 4.900 47.800 ;
        RECT 3.000 47.400 4.900 47.700 ;
        RECT 1.500 45.800 1.800 47.300 ;
        RECT 1.200 45.400 1.800 45.800 ;
        RECT 1.500 45.100 1.800 45.400 ;
        RECT 3.000 45.700 3.400 47.400 ;
        RECT 6.500 47.100 6.900 47.200 ;
        RECT 8.600 47.100 9.000 47.200 ;
        RECT 9.400 47.100 9.700 48.200 ;
        RECT 11.800 47.500 12.200 49.900 ;
        RECT 13.400 48.900 13.800 49.900 ;
        RECT 13.400 47.200 13.700 48.900 ;
        RECT 14.200 47.800 14.600 48.600 ;
        RECT 15.000 47.500 15.400 49.900 ;
        RECT 17.200 49.200 17.600 49.900 ;
        RECT 16.600 48.900 17.600 49.200 ;
        RECT 19.400 48.900 19.800 49.900 ;
        RECT 21.500 49.200 22.100 49.900 ;
        RECT 21.400 48.900 22.100 49.200 ;
        RECT 16.600 48.500 17.000 48.900 ;
        RECT 19.400 48.600 19.700 48.900 ;
        RECT 17.400 48.200 17.800 48.600 ;
        RECT 18.300 48.300 19.700 48.600 ;
        RECT 21.400 48.500 21.800 48.900 ;
        RECT 18.300 48.200 18.700 48.300 ;
        RECT 11.000 47.100 11.800 47.200 ;
        RECT 6.300 46.800 11.800 47.100 ;
        RECT 13.400 46.800 13.800 47.200 ;
        RECT 15.400 47.100 16.200 47.200 ;
        RECT 17.500 47.100 17.800 48.200 ;
        RECT 22.300 47.700 22.700 47.800 ;
        RECT 23.800 47.700 24.200 49.900 ;
        RECT 22.300 47.400 24.200 47.700 ;
        RECT 24.600 47.500 25.000 49.900 ;
        RECT 26.800 49.200 27.200 49.900 ;
        RECT 26.200 48.900 27.200 49.200 ;
        RECT 29.000 48.900 29.400 49.900 ;
        RECT 31.100 49.200 31.700 49.900 ;
        RECT 31.000 48.900 31.700 49.200 ;
        RECT 26.200 48.500 26.600 48.900 ;
        RECT 29.000 48.600 29.300 48.900 ;
        RECT 27.000 47.800 27.400 48.600 ;
        RECT 27.900 48.300 29.300 48.600 ;
        RECT 31.000 48.500 31.400 48.900 ;
        RECT 27.900 48.200 28.300 48.300 ;
        RECT 20.300 47.100 21.000 47.200 ;
        RECT 15.400 46.800 21.000 47.100 ;
        RECT 5.400 46.400 5.800 46.500 ;
        RECT 3.900 46.100 5.800 46.400 ;
        RECT 3.900 46.000 4.300 46.100 ;
        RECT 4.700 45.700 5.100 45.800 ;
        RECT 3.000 45.400 5.100 45.700 ;
        RECT 1.500 44.800 2.600 45.100 ;
        RECT 2.200 41.100 2.600 44.800 ;
        RECT 3.000 41.100 3.400 45.400 ;
        RECT 6.300 45.200 6.600 46.800 ;
        RECT 9.900 46.700 10.300 46.800 ;
        RECT 9.400 46.200 9.800 46.300 ;
        RECT 10.700 46.200 11.100 46.300 ;
        RECT 8.600 45.900 11.100 46.200 ;
        RECT 8.600 45.800 9.000 45.900 ;
        RECT 9.400 45.500 12.200 45.600 ;
        RECT 9.300 45.400 12.200 45.500 ;
        RECT 12.600 45.400 13.000 46.200 ;
        RECT 13.400 46.100 13.700 46.800 ;
        RECT 16.900 46.700 17.300 46.800 ;
        RECT 16.100 46.200 16.500 46.300 ;
        RECT 14.200 46.100 14.600 46.200 ;
        RECT 13.400 45.800 14.600 46.100 ;
        RECT 16.100 45.900 18.600 46.200 ;
        RECT 18.200 45.800 18.600 45.900 ;
        RECT 5.400 44.900 6.600 45.200 ;
        RECT 7.300 45.300 12.200 45.400 ;
        RECT 7.300 45.100 9.700 45.300 ;
        RECT 5.400 44.400 5.700 44.900 ;
        RECT 5.000 44.000 5.700 44.400 ;
        RECT 6.500 44.500 6.900 44.600 ;
        RECT 7.300 44.500 7.600 45.100 ;
        RECT 6.500 44.200 7.600 44.500 ;
        RECT 7.900 44.500 10.600 44.800 ;
        RECT 7.900 44.400 8.300 44.500 ;
        RECT 10.200 44.400 10.600 44.500 ;
        RECT 7.100 43.700 7.500 43.800 ;
        RECT 8.500 43.700 8.900 43.800 ;
        RECT 5.400 43.100 5.800 43.500 ;
        RECT 7.100 43.400 8.900 43.700 ;
        RECT 7.500 43.100 7.800 43.400 ;
        RECT 10.200 43.100 10.600 43.500 ;
        RECT 5.100 41.100 5.700 43.100 ;
        RECT 7.400 41.100 7.800 43.100 ;
        RECT 9.600 42.800 10.600 43.100 ;
        RECT 9.600 41.100 10.000 42.800 ;
        RECT 11.800 41.100 12.200 45.300 ;
        RECT 13.400 45.100 13.700 45.800 ;
        RECT 15.000 45.500 17.800 45.600 ;
        RECT 15.000 45.400 17.900 45.500 ;
        RECT 15.000 45.300 19.900 45.400 ;
        RECT 12.900 44.700 13.800 45.100 ;
        RECT 12.900 41.100 13.300 44.700 ;
        RECT 15.000 41.100 15.400 45.300 ;
        RECT 17.500 45.100 19.900 45.300 ;
        RECT 16.600 44.500 19.300 44.800 ;
        RECT 16.600 44.400 17.000 44.500 ;
        RECT 18.900 44.400 19.300 44.500 ;
        RECT 19.600 44.500 19.900 45.100 ;
        RECT 20.600 45.200 20.900 46.800 ;
        RECT 21.400 46.400 21.800 46.500 ;
        RECT 21.400 46.100 23.300 46.400 ;
        RECT 22.900 46.000 23.300 46.100 ;
        RECT 22.100 45.700 22.500 45.800 ;
        RECT 23.800 45.700 24.200 47.400 ;
        RECT 25.000 47.100 25.800 47.200 ;
        RECT 27.100 47.100 27.400 47.800 ;
        RECT 31.900 47.700 32.300 47.800 ;
        RECT 33.400 47.700 33.800 49.900 ;
        RECT 36.600 48.900 37.000 49.900 ;
        RECT 38.200 49.200 38.600 49.900 ;
        RECT 31.900 47.400 33.800 47.700 ;
        RECT 29.900 47.100 30.300 47.200 ;
        RECT 25.000 46.800 30.500 47.100 ;
        RECT 26.500 46.700 26.900 46.800 ;
        RECT 25.700 46.200 26.100 46.300 ;
        RECT 30.200 46.200 30.500 46.800 ;
        RECT 31.000 46.400 31.400 46.500 ;
        RECT 25.700 45.900 28.200 46.200 ;
        RECT 27.800 45.800 28.200 45.900 ;
        RECT 30.200 45.800 30.600 46.200 ;
        RECT 31.000 46.100 32.900 46.400 ;
        RECT 32.500 46.000 32.900 46.100 ;
        RECT 22.100 45.400 24.200 45.700 ;
        RECT 20.600 44.900 21.800 45.200 ;
        RECT 20.300 44.500 20.700 44.600 ;
        RECT 19.600 44.200 20.700 44.500 ;
        RECT 21.500 44.400 21.800 44.900 ;
        RECT 21.500 44.000 22.200 44.400 ;
        RECT 18.300 43.700 18.700 43.800 ;
        RECT 19.700 43.700 20.100 43.800 ;
        RECT 16.600 43.100 17.000 43.500 ;
        RECT 18.300 43.400 20.100 43.700 ;
        RECT 19.400 43.100 19.700 43.400 ;
        RECT 21.400 43.100 21.800 43.500 ;
        RECT 16.600 42.800 17.600 43.100 ;
        RECT 17.200 41.100 17.600 42.800 ;
        RECT 19.400 41.100 19.800 43.100 ;
        RECT 21.500 41.100 22.100 43.100 ;
        RECT 23.800 41.100 24.200 45.400 ;
        RECT 24.600 45.500 27.400 45.600 ;
        RECT 24.600 45.400 27.500 45.500 ;
        RECT 24.600 45.300 29.500 45.400 ;
        RECT 24.600 41.100 25.000 45.300 ;
        RECT 27.100 45.100 29.500 45.300 ;
        RECT 26.200 44.500 28.900 44.800 ;
        RECT 26.200 44.400 26.600 44.500 ;
        RECT 28.500 44.400 28.900 44.500 ;
        RECT 29.200 44.500 29.500 45.100 ;
        RECT 30.200 45.200 30.500 45.800 ;
        RECT 31.700 45.700 32.100 45.800 ;
        RECT 33.400 45.700 33.800 47.400 ;
        RECT 31.700 45.400 33.800 45.700 ;
        RECT 30.200 44.900 31.400 45.200 ;
        RECT 29.900 44.500 30.300 44.600 ;
        RECT 29.200 44.200 30.300 44.500 ;
        RECT 31.100 44.400 31.400 44.900 ;
        RECT 31.100 44.000 31.800 44.400 ;
        RECT 27.900 43.700 28.300 43.800 ;
        RECT 29.300 43.700 29.700 43.800 ;
        RECT 26.200 43.100 26.600 43.500 ;
        RECT 27.900 43.400 29.700 43.700 ;
        RECT 29.000 43.100 29.300 43.400 ;
        RECT 31.000 43.100 31.400 43.500 ;
        RECT 26.200 42.800 27.200 43.100 ;
        RECT 26.800 41.100 27.200 42.800 ;
        RECT 29.000 41.100 29.400 43.100 ;
        RECT 31.100 41.100 31.700 43.100 ;
        RECT 33.400 41.100 33.800 45.400 ;
        RECT 36.400 48.800 37.000 48.900 ;
        RECT 38.100 48.800 38.600 49.200 ;
        RECT 36.400 48.500 38.400 48.800 ;
        RECT 36.400 45.200 36.700 48.500 ;
        RECT 38.500 47.800 39.400 48.200 ;
        RECT 40.600 47.900 41.000 49.900 ;
        RECT 42.800 49.200 43.600 49.900 ;
        RECT 42.200 48.800 43.600 49.200 ;
        RECT 42.800 48.100 43.600 48.800 ;
        RECT 40.600 47.600 41.800 47.900 ;
        RECT 41.400 47.500 41.800 47.600 ;
        RECT 42.100 47.400 42.500 47.800 ;
        RECT 42.100 47.200 42.400 47.400 ;
        RECT 37.800 46.800 38.600 47.200 ;
        RECT 40.600 46.800 41.400 47.200 ;
        RECT 42.000 46.800 42.400 47.200 ;
        RECT 42.800 47.100 43.100 48.100 ;
        RECT 45.400 47.900 45.800 49.900 ;
        RECT 43.400 47.400 44.200 47.800 ;
        RECT 44.500 47.600 45.800 47.900 ;
        RECT 47.800 47.700 48.200 49.900 ;
        RECT 49.900 49.200 50.500 49.900 ;
        RECT 49.900 48.900 50.600 49.200 ;
        RECT 52.200 48.900 52.600 49.900 ;
        RECT 54.400 49.200 54.800 49.900 ;
        RECT 54.400 48.900 55.400 49.200 ;
        RECT 50.200 48.500 50.600 48.900 ;
        RECT 52.300 48.600 52.600 48.900 ;
        RECT 52.300 48.300 53.700 48.600 ;
        RECT 53.300 48.200 53.700 48.300 ;
        RECT 54.200 48.200 54.600 48.600 ;
        RECT 55.000 48.500 55.400 48.900 ;
        RECT 49.300 47.700 49.700 47.800 ;
        RECT 44.500 47.500 44.900 47.600 ;
        RECT 47.800 47.400 49.700 47.700 ;
        RECT 45.000 47.100 45.800 47.200 ;
        RECT 42.800 46.800 43.300 47.100 ;
        RECT 44.700 47.000 45.800 47.100 ;
        RECT 43.000 46.200 43.300 46.800 ;
        RECT 43.600 46.800 45.800 47.000 ;
        RECT 43.600 46.700 45.000 46.800 ;
        RECT 43.600 46.600 44.000 46.700 ;
        RECT 37.000 46.100 37.800 46.200 ;
        RECT 42.200 46.100 42.600 46.200 ;
        RECT 37.000 45.800 42.600 46.100 ;
        RECT 43.000 45.800 43.400 46.200 ;
        RECT 44.300 46.100 44.700 46.200 ;
        RECT 43.900 45.800 44.700 46.100 ;
        RECT 35.000 44.900 36.700 45.200 ;
        RECT 43.000 45.100 43.300 45.800 ;
        RECT 43.900 45.700 44.300 45.800 ;
        RECT 47.800 45.700 48.200 47.400 ;
        RECT 51.300 47.100 51.700 47.200 ;
        RECT 54.200 47.100 54.500 48.200 ;
        RECT 56.600 47.500 57.000 49.900 ;
        RECT 58.200 47.600 58.600 49.900 ;
        RECT 59.800 47.600 60.200 49.900 ;
        RECT 61.400 47.600 61.800 49.900 ;
        RECT 63.000 47.600 63.400 49.900 ;
        RECT 57.400 47.200 58.600 47.600 ;
        RECT 59.100 47.200 60.200 47.600 ;
        RECT 60.700 47.200 61.800 47.600 ;
        RECT 62.500 47.200 63.400 47.600 ;
        RECT 55.800 47.100 56.600 47.200 ;
        RECT 51.100 46.800 56.600 47.100 ;
        RECT 50.200 46.400 50.600 46.500 ;
        RECT 48.700 46.100 50.600 46.400 ;
        RECT 48.700 46.000 49.100 46.100 ;
        RECT 49.500 45.700 49.900 45.800 ;
        RECT 47.800 45.400 49.900 45.700 ;
        RECT 35.000 44.800 35.400 44.900 ;
        RECT 35.100 44.500 35.400 44.800 ;
        RECT 40.600 44.800 41.800 45.100 ;
        RECT 35.900 44.500 37.700 44.600 ;
        RECT 34.200 41.500 34.600 44.500 ;
        RECT 35.000 41.700 35.400 44.500 ;
        RECT 35.800 44.300 37.700 44.500 ;
        RECT 34.300 41.400 34.600 41.500 ;
        RECT 35.800 41.500 36.200 44.300 ;
        RECT 37.400 44.100 37.700 44.300 ;
        RECT 38.300 44.400 40.100 44.700 ;
        RECT 38.300 44.100 38.600 44.400 ;
        RECT 35.800 41.400 36.100 41.500 ;
        RECT 34.300 41.100 36.100 41.400 ;
        RECT 36.600 41.400 37.000 44.000 ;
        RECT 37.400 41.700 37.800 44.100 ;
        RECT 38.200 41.400 38.600 44.100 ;
        RECT 36.600 41.100 38.600 41.400 ;
        RECT 39.800 44.100 40.100 44.400 ;
        RECT 39.800 41.100 40.200 44.100 ;
        RECT 40.600 41.100 41.000 44.800 ;
        RECT 41.400 44.700 41.800 44.800 ;
        RECT 42.800 41.100 43.600 45.100 ;
        RECT 44.500 44.800 45.800 45.100 ;
        RECT 44.500 44.700 44.900 44.800 ;
        RECT 45.400 41.100 45.800 44.800 ;
        RECT 47.800 41.100 48.200 45.400 ;
        RECT 51.100 45.200 51.400 46.800 ;
        RECT 54.700 46.700 55.100 46.800 ;
        RECT 54.200 46.200 54.600 46.300 ;
        RECT 55.500 46.200 55.900 46.300 ;
        RECT 53.400 45.900 55.900 46.200 ;
        RECT 53.400 45.800 53.800 45.900 ;
        RECT 57.400 45.800 57.800 47.200 ;
        RECT 59.100 46.900 59.500 47.200 ;
        RECT 60.700 46.900 61.100 47.200 ;
        RECT 62.500 46.900 62.900 47.200 ;
        RECT 58.200 46.500 59.500 46.900 ;
        RECT 59.900 46.500 61.100 46.900 ;
        RECT 61.600 46.500 62.900 46.900 ;
        RECT 59.100 45.800 59.500 46.500 ;
        RECT 60.700 45.800 61.100 46.500 ;
        RECT 62.500 45.800 62.900 46.500 ;
        RECT 64.600 46.200 65.000 49.900 ;
        RECT 66.200 47.600 66.600 49.900 ;
        RECT 65.500 47.300 66.600 47.600 ;
        RECT 54.200 45.500 57.000 45.600 ;
        RECT 54.100 45.400 57.000 45.500 ;
        RECT 57.400 45.400 58.600 45.800 ;
        RECT 59.100 45.400 60.200 45.800 ;
        RECT 60.700 45.400 61.800 45.800 ;
        RECT 62.500 45.400 63.400 45.800 ;
        RECT 50.200 44.900 51.400 45.200 ;
        RECT 52.100 45.300 57.000 45.400 ;
        RECT 52.100 45.100 54.500 45.300 ;
        RECT 50.200 44.400 50.500 44.900 ;
        RECT 49.800 44.000 50.500 44.400 ;
        RECT 51.300 44.500 51.700 44.600 ;
        RECT 52.100 44.500 52.400 45.100 ;
        RECT 51.300 44.200 52.400 44.500 ;
        RECT 52.700 44.500 55.400 44.800 ;
        RECT 52.700 44.400 53.100 44.500 ;
        RECT 55.000 44.400 55.400 44.500 ;
        RECT 51.900 43.700 52.300 43.800 ;
        RECT 53.300 43.700 53.700 43.800 ;
        RECT 50.200 43.100 50.600 43.500 ;
        RECT 51.900 43.400 53.700 43.700 ;
        RECT 52.300 43.100 52.600 43.400 ;
        RECT 55.000 43.100 55.400 43.500 ;
        RECT 49.900 41.100 50.500 43.100 ;
        RECT 52.200 41.100 52.600 43.100 ;
        RECT 54.400 42.800 55.400 43.100 ;
        RECT 54.400 41.100 54.800 42.800 ;
        RECT 56.600 41.100 57.000 45.300 ;
        RECT 58.200 41.100 58.600 45.400 ;
        RECT 59.800 41.100 60.200 45.400 ;
        RECT 61.400 41.100 61.800 45.400 ;
        RECT 63.000 41.100 63.400 45.400 ;
        RECT 64.600 45.100 64.900 46.200 ;
        RECT 65.500 45.800 65.800 47.300 ;
        RECT 66.200 46.100 66.600 46.600 ;
        RECT 67.000 46.100 67.400 49.900 ;
        RECT 67.800 47.800 68.200 48.600 ;
        RECT 66.200 45.800 67.400 46.100 ;
        RECT 65.200 45.400 65.800 45.800 ;
        RECT 65.500 45.100 65.800 45.400 ;
        RECT 64.600 41.100 65.000 45.100 ;
        RECT 65.500 44.800 66.600 45.100 ;
        RECT 66.200 41.100 66.600 44.800 ;
        RECT 67.000 41.100 67.400 45.800 ;
        RECT 68.600 47.700 69.000 49.900 ;
        RECT 70.700 49.200 71.300 49.900 ;
        RECT 70.700 48.900 71.400 49.200 ;
        RECT 73.000 48.900 73.400 49.900 ;
        RECT 75.200 49.200 75.600 49.900 ;
        RECT 75.200 48.900 76.200 49.200 ;
        RECT 71.000 48.500 71.400 48.900 ;
        RECT 73.100 48.600 73.400 48.900 ;
        RECT 73.100 48.300 74.500 48.600 ;
        RECT 74.100 48.200 74.500 48.300 ;
        RECT 75.000 48.200 75.400 48.600 ;
        RECT 75.800 48.500 76.200 48.900 ;
        RECT 70.100 47.700 70.500 47.800 ;
        RECT 68.600 47.400 70.500 47.700 ;
        RECT 68.600 45.700 69.000 47.400 ;
        RECT 72.100 47.100 72.500 47.200 ;
        RECT 73.400 47.100 73.800 47.200 ;
        RECT 75.000 47.100 75.300 48.200 ;
        RECT 77.400 47.500 77.800 49.900 ;
        RECT 78.200 47.900 78.600 49.900 ;
        RECT 79.000 48.000 79.400 49.900 ;
        RECT 80.600 48.000 81.000 49.900 ;
        RECT 82.700 48.200 83.100 49.900 ;
        RECT 79.000 47.900 81.000 48.000 ;
        RECT 82.200 47.900 83.100 48.200 ;
        RECT 84.600 48.900 85.000 49.900 ;
        RECT 78.300 47.200 78.600 47.900 ;
        RECT 79.100 47.700 80.900 47.900 ;
        RECT 80.200 47.200 80.600 47.400 ;
        RECT 76.600 47.100 77.400 47.200 ;
        RECT 71.900 46.800 77.400 47.100 ;
        RECT 78.200 46.800 79.500 47.200 ;
        RECT 80.200 46.900 81.000 47.200 ;
        RECT 80.600 46.800 81.000 46.900 ;
        RECT 81.400 46.800 81.800 47.600 ;
        RECT 71.000 46.400 71.400 46.500 ;
        RECT 69.500 46.100 71.400 46.400 ;
        RECT 69.500 46.000 69.900 46.100 ;
        RECT 70.300 45.700 70.700 45.800 ;
        RECT 68.600 45.400 70.700 45.700 ;
        RECT 68.600 41.100 69.000 45.400 ;
        RECT 71.900 45.200 72.200 46.800 ;
        RECT 75.500 46.700 75.900 46.800 ;
        RECT 76.300 46.200 76.700 46.300 ;
        RECT 74.200 45.900 76.700 46.200 ;
        RECT 74.200 45.800 74.600 45.900 ;
        RECT 75.000 45.500 77.800 45.600 ;
        RECT 74.900 45.400 77.800 45.500 ;
        RECT 71.000 44.900 72.200 45.200 ;
        RECT 72.900 45.300 77.800 45.400 ;
        RECT 72.900 45.100 75.300 45.300 ;
        RECT 71.000 44.400 71.300 44.900 ;
        RECT 70.600 44.000 71.300 44.400 ;
        RECT 72.100 44.500 72.500 44.600 ;
        RECT 72.900 44.500 73.200 45.100 ;
        RECT 72.100 44.200 73.200 44.500 ;
        RECT 73.500 44.500 76.200 44.800 ;
        RECT 73.500 44.400 73.900 44.500 ;
        RECT 75.800 44.400 76.200 44.500 ;
        RECT 72.700 43.700 73.100 43.800 ;
        RECT 74.100 43.700 74.500 43.800 ;
        RECT 71.000 43.100 71.400 43.500 ;
        RECT 72.700 43.400 74.500 43.700 ;
        RECT 73.100 43.100 73.400 43.400 ;
        RECT 75.800 43.100 76.200 43.500 ;
        RECT 70.700 41.100 71.300 43.100 ;
        RECT 73.000 41.100 73.400 43.100 ;
        RECT 75.200 42.800 76.200 43.100 ;
        RECT 75.200 41.100 75.600 42.800 ;
        RECT 77.400 41.100 77.800 45.300 ;
        RECT 78.200 45.100 78.600 45.200 ;
        RECT 79.200 45.100 79.500 46.800 ;
        RECT 79.800 46.100 80.200 46.600 ;
        RECT 81.400 46.100 81.700 46.800 ;
        RECT 79.800 45.800 81.700 46.100 ;
        RECT 82.200 46.100 82.600 47.900 ;
        RECT 84.600 47.200 84.900 48.900 ;
        RECT 85.400 48.100 85.800 48.600 ;
        RECT 86.200 48.100 86.600 49.900 ;
        RECT 88.600 48.800 89.000 49.900 ;
        RECT 85.400 47.800 86.600 48.100 ;
        RECT 84.600 46.800 85.000 47.200 ;
        RECT 83.800 46.100 84.200 46.200 ;
        RECT 82.200 45.800 84.200 46.100 ;
        RECT 78.200 44.800 78.900 45.100 ;
        RECT 79.200 44.800 79.700 45.100 ;
        RECT 78.600 44.200 78.900 44.800 ;
        RECT 78.600 43.800 79.000 44.200 ;
        RECT 79.300 41.100 79.700 44.800 ;
        RECT 82.200 41.100 82.600 45.800 ;
        RECT 83.800 45.400 84.200 45.800 ;
        RECT 84.600 45.200 84.900 46.800 ;
        RECT 83.000 44.400 83.400 45.200 ;
        RECT 84.600 45.100 85.000 45.200 ;
        RECT 84.100 44.700 85.000 45.100 ;
        RECT 84.100 41.100 84.500 44.700 ;
        RECT 86.200 41.100 86.600 47.800 ;
        RECT 87.800 47.800 88.200 48.600 ;
        RECT 87.000 47.100 87.400 47.600 ;
        RECT 87.800 47.200 88.100 47.800 ;
        RECT 88.700 47.200 89.000 48.800 ;
        RECT 91.500 48.200 91.900 49.900 ;
        RECT 91.000 47.900 91.900 48.200 ;
        RECT 87.800 47.100 88.200 47.200 ;
        RECT 87.000 46.800 88.200 47.100 ;
        RECT 88.600 46.800 89.000 47.200 ;
        RECT 90.200 46.800 90.600 47.600 ;
        RECT 88.700 45.100 89.000 46.800 ;
        RECT 89.400 46.100 89.800 46.200 ;
        RECT 91.000 46.100 91.400 47.900 ;
        RECT 92.600 46.800 93.000 47.600 ;
        RECT 89.400 45.800 91.400 46.100 ;
        RECT 89.400 45.400 89.800 45.800 ;
        RECT 90.200 45.100 90.600 45.200 ;
        RECT 91.000 45.100 91.400 45.800 ;
        RECT 88.600 44.700 89.500 45.100 ;
        RECT 90.200 44.800 91.400 45.100 ;
        RECT 89.100 41.100 89.500 44.700 ;
        RECT 91.000 41.100 91.400 44.800 ;
        RECT 91.800 44.400 92.200 45.200 ;
        RECT 93.400 41.100 93.800 49.900 ;
        RECT 98.200 48.900 98.600 49.900 ;
        RECT 99.800 49.200 100.200 49.900 ;
        RECT 98.000 48.800 98.600 48.900 ;
        RECT 99.700 48.800 100.200 49.200 ;
        RECT 98.000 48.500 100.000 48.800 ;
        RECT 98.000 45.200 98.300 48.500 ;
        RECT 99.800 47.800 101.000 48.200 ;
        RECT 99.400 47.100 100.200 47.200 ;
        RECT 102.200 47.100 102.600 49.900 ;
        RECT 103.000 47.800 103.400 48.600 ;
        RECT 103.800 47.600 104.200 49.900 ;
        RECT 103.800 47.300 104.900 47.600 ;
        RECT 99.400 46.800 102.600 47.100 ;
        RECT 98.600 45.800 99.400 46.200 ;
        RECT 96.600 44.900 98.300 45.200 ;
        RECT 96.600 44.800 97.000 44.900 ;
        RECT 96.700 44.500 97.000 44.800 ;
        RECT 97.500 44.500 99.300 44.600 ;
        RECT 95.800 41.500 96.200 44.500 ;
        RECT 96.600 41.700 97.000 44.500 ;
        RECT 97.400 44.300 99.300 44.500 ;
        RECT 95.900 41.400 96.200 41.500 ;
        RECT 97.400 41.500 97.800 44.300 ;
        RECT 99.000 44.100 99.300 44.300 ;
        RECT 99.900 44.400 101.700 44.700 ;
        RECT 99.900 44.100 100.200 44.400 ;
        RECT 97.400 41.400 97.700 41.500 ;
        RECT 95.900 41.100 97.700 41.400 ;
        RECT 98.200 41.400 98.600 44.000 ;
        RECT 99.000 41.700 99.400 44.100 ;
        RECT 99.800 41.400 100.200 44.100 ;
        RECT 98.200 41.100 100.200 41.400 ;
        RECT 101.400 44.100 101.700 44.400 ;
        RECT 101.400 41.100 101.800 44.100 ;
        RECT 102.200 41.100 102.600 46.800 ;
        RECT 103.000 46.100 103.400 46.200 ;
        RECT 103.800 46.100 104.200 46.600 ;
        RECT 103.000 45.800 104.200 46.100 ;
        RECT 104.600 45.800 104.900 47.300 ;
        RECT 105.400 46.200 105.800 49.900 ;
        RECT 107.800 49.200 108.200 49.900 ;
        RECT 107.800 48.900 108.300 49.200 ;
        RECT 108.000 48.800 108.300 48.900 ;
        RECT 109.400 49.100 109.800 49.900 ;
        RECT 114.100 49.200 114.900 49.900 ;
        RECT 111.800 49.100 112.200 49.200 ;
        RECT 109.400 48.800 112.200 49.100 ;
        RECT 114.100 48.800 115.400 49.200 ;
        RECT 108.000 48.500 110.000 48.800 ;
        RECT 107.000 47.800 107.900 48.200 ;
        RECT 107.800 46.800 108.600 47.200 ;
        RECT 104.600 45.400 105.200 45.800 ;
        RECT 104.600 45.100 104.900 45.400 ;
        RECT 105.500 45.100 105.800 46.200 ;
        RECT 108.600 45.800 109.400 46.200 ;
        RECT 103.800 44.800 104.900 45.100 ;
        RECT 103.800 41.100 104.200 44.800 ;
        RECT 105.400 41.100 105.800 45.100 ;
        RECT 109.700 45.200 110.000 48.500 ;
        RECT 114.100 47.900 114.900 48.800 ;
        RECT 118.200 47.900 118.600 49.900 ;
        RECT 118.900 48.200 119.300 48.600 ;
        RECT 113.400 46.400 113.800 47.200 ;
        RECT 114.300 46.200 114.600 47.900 ;
        RECT 115.000 46.800 115.400 47.200 ;
        RECT 117.400 47.100 117.800 47.200 ;
        RECT 115.800 46.800 117.800 47.100 ;
        RECT 115.000 46.600 115.300 46.800 ;
        RECT 114.900 46.200 115.300 46.600 ;
        RECT 115.800 46.200 116.100 46.800 ;
        RECT 117.400 46.400 117.800 46.800 ;
        RECT 112.600 46.100 113.000 46.200 ;
        RECT 112.600 45.800 113.400 46.100 ;
        RECT 114.200 45.800 114.600 46.200 ;
        RECT 113.000 45.600 113.400 45.800 ;
        RECT 114.300 45.700 114.600 45.800 ;
        RECT 114.300 45.400 115.300 45.700 ;
        RECT 115.800 45.400 116.200 46.200 ;
        RECT 116.600 46.100 117.000 46.200 ;
        RECT 118.200 46.100 118.500 47.900 ;
        RECT 119.000 47.800 119.400 48.200 ;
        RECT 119.800 47.700 120.200 49.900 ;
        RECT 121.900 49.200 122.500 49.900 ;
        RECT 121.900 48.900 122.600 49.200 ;
        RECT 124.200 48.900 124.600 49.900 ;
        RECT 126.400 49.200 126.800 49.900 ;
        RECT 126.400 48.900 127.400 49.200 ;
        RECT 122.200 48.500 122.600 48.900 ;
        RECT 124.300 48.600 124.600 48.900 ;
        RECT 124.300 48.300 125.700 48.600 ;
        RECT 125.300 48.200 125.700 48.300 ;
        RECT 126.200 48.200 126.600 48.600 ;
        RECT 127.000 48.500 127.400 48.900 ;
        RECT 121.300 47.700 121.700 47.800 ;
        RECT 119.800 47.400 121.700 47.700 ;
        RECT 119.000 46.100 119.400 46.200 ;
        RECT 116.600 45.800 117.400 46.100 ;
        RECT 118.200 45.800 119.400 46.100 ;
        RECT 117.000 45.600 117.400 45.800 ;
        RECT 109.700 44.900 111.400 45.200 ;
        RECT 115.000 45.100 115.300 45.400 ;
        RECT 119.000 45.100 119.300 45.800 ;
        RECT 119.800 45.700 120.200 47.400 ;
        RECT 123.300 47.100 123.700 47.200 ;
        RECT 126.200 47.100 126.500 48.200 ;
        RECT 128.600 47.500 129.000 49.900 ;
        RECT 129.400 47.500 129.800 49.900 ;
        RECT 131.600 49.200 132.000 49.900 ;
        RECT 131.000 48.900 132.000 49.200 ;
        RECT 133.800 48.900 134.200 49.900 ;
        RECT 135.900 49.200 136.500 49.900 ;
        RECT 135.800 48.900 136.500 49.200 ;
        RECT 138.200 49.100 138.600 49.900 ;
        RECT 139.000 49.100 139.400 49.900 ;
        RECT 131.000 48.500 131.400 48.900 ;
        RECT 133.800 48.600 134.100 48.900 ;
        RECT 131.800 48.200 132.200 48.600 ;
        RECT 132.700 48.300 134.100 48.600 ;
        RECT 135.800 48.500 136.200 48.900 ;
        RECT 138.200 48.800 139.400 49.100 ;
        RECT 141.100 49.200 141.700 49.900 ;
        RECT 141.100 48.900 141.800 49.200 ;
        RECT 143.400 48.900 143.800 49.900 ;
        RECT 145.600 49.200 146.000 49.900 ;
        RECT 145.600 48.900 146.600 49.200 ;
        RECT 132.700 48.200 133.100 48.300 ;
        RECT 127.800 47.100 128.600 47.200 ;
        RECT 129.800 47.100 130.600 47.200 ;
        RECT 131.900 47.100 132.200 48.200 ;
        RECT 136.700 47.700 137.100 47.800 ;
        RECT 138.200 47.700 138.600 48.800 ;
        RECT 136.700 47.400 138.600 47.700 ;
        RECT 134.700 47.100 135.100 47.200 ;
        RECT 123.100 46.800 135.300 47.100 ;
        RECT 122.200 46.400 122.600 46.500 ;
        RECT 120.700 46.100 122.600 46.400 ;
        RECT 120.700 46.000 121.100 46.100 ;
        RECT 121.500 45.700 121.900 45.800 ;
        RECT 119.800 45.400 121.900 45.700 ;
        RECT 111.000 44.800 111.400 44.900 ;
        RECT 112.600 44.800 114.600 45.100 ;
        RECT 106.300 44.400 108.100 44.700 ;
        RECT 106.300 44.100 106.600 44.400 ;
        RECT 106.200 41.100 106.600 44.100 ;
        RECT 107.800 44.100 108.100 44.400 ;
        RECT 108.700 44.500 110.500 44.600 ;
        RECT 111.000 44.500 111.300 44.800 ;
        RECT 108.700 44.300 110.600 44.500 ;
        RECT 108.700 44.100 109.000 44.300 ;
        RECT 107.800 41.400 108.200 44.100 ;
        RECT 108.600 41.700 109.000 44.100 ;
        RECT 109.400 41.400 109.800 44.000 ;
        RECT 110.200 41.500 110.600 44.300 ;
        RECT 111.000 41.700 111.400 44.500 ;
        RECT 107.800 41.100 109.800 41.400 ;
        RECT 110.300 41.400 110.600 41.500 ;
        RECT 111.800 41.500 112.200 44.500 ;
        RECT 111.800 41.400 112.100 41.500 ;
        RECT 110.300 41.100 112.100 41.400 ;
        RECT 112.600 41.100 113.000 44.800 ;
        RECT 114.200 41.400 114.600 44.800 ;
        RECT 115.000 41.700 115.400 45.100 ;
        RECT 115.800 41.400 116.200 45.100 ;
        RECT 114.200 41.100 116.200 41.400 ;
        RECT 116.600 44.800 118.600 45.100 ;
        RECT 116.600 41.100 117.000 44.800 ;
        RECT 118.200 41.100 118.600 44.800 ;
        RECT 119.000 41.100 119.400 45.100 ;
        RECT 119.800 41.100 120.200 45.400 ;
        RECT 123.100 45.200 123.400 46.800 ;
        RECT 126.700 46.700 127.100 46.800 ;
        RECT 131.300 46.700 131.700 46.800 ;
        RECT 126.200 46.200 126.600 46.300 ;
        RECT 127.500 46.200 127.900 46.300 ;
        RECT 125.400 45.900 127.900 46.200 ;
        RECT 130.500 46.200 130.900 46.300 ;
        RECT 130.500 45.900 133.000 46.200 ;
        RECT 125.400 45.800 125.800 45.900 ;
        RECT 132.600 45.800 133.000 45.900 ;
        RECT 126.200 45.500 129.000 45.600 ;
        RECT 126.100 45.400 129.000 45.500 ;
        RECT 122.200 44.900 123.400 45.200 ;
        RECT 124.100 45.300 129.000 45.400 ;
        RECT 124.100 45.100 126.500 45.300 ;
        RECT 122.200 44.400 122.500 44.900 ;
        RECT 121.800 44.200 122.500 44.400 ;
        RECT 123.300 44.500 123.700 44.600 ;
        RECT 124.100 44.500 124.400 45.100 ;
        RECT 123.300 44.200 124.400 44.500 ;
        RECT 124.700 44.500 127.400 44.800 ;
        RECT 124.700 44.400 125.100 44.500 ;
        RECT 127.000 44.400 127.400 44.500 ;
        RECT 121.400 44.000 122.500 44.200 ;
        RECT 121.400 43.800 122.100 44.000 ;
        RECT 123.900 43.700 124.300 43.800 ;
        RECT 125.300 43.700 125.700 43.800 ;
        RECT 122.200 43.100 122.600 43.500 ;
        RECT 123.900 43.400 125.700 43.700 ;
        RECT 124.300 43.100 124.600 43.400 ;
        RECT 127.000 43.100 127.400 43.500 ;
        RECT 121.900 41.100 122.500 43.100 ;
        RECT 124.200 41.100 124.600 43.100 ;
        RECT 126.400 42.800 127.400 43.100 ;
        RECT 126.400 41.100 126.800 42.800 ;
        RECT 128.600 41.100 129.000 45.300 ;
        RECT 129.400 45.500 132.200 45.600 ;
        RECT 129.400 45.400 132.300 45.500 ;
        RECT 129.400 45.300 134.300 45.400 ;
        RECT 129.400 41.100 129.800 45.300 ;
        RECT 131.900 45.100 134.300 45.300 ;
        RECT 131.000 44.500 133.700 44.800 ;
        RECT 131.000 44.400 131.400 44.500 ;
        RECT 133.300 44.400 133.700 44.500 ;
        RECT 134.000 44.500 134.300 45.100 ;
        RECT 135.000 45.200 135.300 46.800 ;
        RECT 135.800 46.400 136.200 46.500 ;
        RECT 135.800 46.100 137.700 46.400 ;
        RECT 137.300 46.000 137.700 46.100 ;
        RECT 136.500 45.700 136.900 45.800 ;
        RECT 138.200 45.700 138.600 47.400 ;
        RECT 136.500 45.400 138.600 45.700 ;
        RECT 135.000 44.900 136.200 45.200 ;
        RECT 134.700 44.500 135.100 44.600 ;
        RECT 134.000 44.200 135.100 44.500 ;
        RECT 135.900 44.400 136.200 44.900 ;
        RECT 135.900 44.000 136.600 44.400 ;
        RECT 132.700 43.700 133.100 43.800 ;
        RECT 134.100 43.700 134.500 43.800 ;
        RECT 131.000 43.100 131.400 43.500 ;
        RECT 132.700 43.400 134.500 43.700 ;
        RECT 133.800 43.100 134.100 43.400 ;
        RECT 135.800 43.100 136.200 43.500 ;
        RECT 131.000 42.800 132.000 43.100 ;
        RECT 131.600 41.100 132.000 42.800 ;
        RECT 133.800 41.100 134.200 43.100 ;
        RECT 135.900 41.100 136.500 43.100 ;
        RECT 138.200 41.100 138.600 45.400 ;
        RECT 139.000 47.700 139.400 48.800 ;
        RECT 141.400 48.500 141.800 48.900 ;
        RECT 143.500 48.600 143.800 48.900 ;
        RECT 143.500 48.300 144.900 48.600 ;
        RECT 144.500 48.200 144.900 48.300 ;
        RECT 145.400 48.200 145.800 48.600 ;
        RECT 146.200 48.500 146.600 48.900 ;
        RECT 140.500 47.700 140.900 47.800 ;
        RECT 139.000 47.400 140.900 47.700 ;
        RECT 139.000 45.700 139.400 47.400 ;
        RECT 142.500 47.100 142.900 47.200 ;
        RECT 144.600 47.100 145.000 47.200 ;
        RECT 145.400 47.100 145.700 48.200 ;
        RECT 147.800 47.500 148.200 49.900 ;
        RECT 151.000 48.900 151.400 49.900 ;
        RECT 153.400 48.900 153.800 49.900 ;
        RECT 150.200 47.800 150.600 48.600 ;
        RECT 151.100 48.200 151.400 48.900 ;
        RECT 151.000 47.800 151.400 48.200 ;
        RECT 152.600 47.800 153.000 48.600 ;
        RECT 151.100 47.200 151.400 47.800 ;
        RECT 153.500 47.200 153.800 48.900 ;
        RECT 147.000 47.100 147.800 47.200 ;
        RECT 142.300 46.800 147.800 47.100 ;
        RECT 151.000 46.800 151.400 47.200 ;
        RECT 141.400 46.400 141.800 46.500 ;
        RECT 139.900 46.100 141.800 46.400 ;
        RECT 139.900 46.000 140.300 46.100 ;
        RECT 140.700 45.700 141.100 45.800 ;
        RECT 139.000 45.400 141.100 45.700 ;
        RECT 139.000 41.100 139.400 45.400 ;
        RECT 142.300 45.200 142.600 46.800 ;
        RECT 145.900 46.700 146.300 46.800 ;
        RECT 145.400 46.200 145.800 46.300 ;
        RECT 146.700 46.200 147.100 46.300 ;
        RECT 144.600 45.900 147.100 46.200 ;
        RECT 144.600 45.800 145.000 45.900 ;
        RECT 145.400 45.500 148.200 45.600 ;
        RECT 145.300 45.400 148.200 45.500 ;
        RECT 141.400 44.900 142.600 45.200 ;
        RECT 143.300 45.300 148.200 45.400 ;
        RECT 143.300 45.100 145.700 45.300 ;
        RECT 141.400 44.400 141.700 44.900 ;
        RECT 141.000 44.000 141.700 44.400 ;
        RECT 142.500 44.500 142.900 44.600 ;
        RECT 143.300 44.500 143.600 45.100 ;
        RECT 142.500 44.200 143.600 44.500 ;
        RECT 143.900 44.500 146.600 44.800 ;
        RECT 143.900 44.400 144.300 44.500 ;
        RECT 146.200 44.400 146.600 44.500 ;
        RECT 143.100 43.700 143.500 43.800 ;
        RECT 144.500 43.700 144.900 43.800 ;
        RECT 141.400 43.100 141.800 43.500 ;
        RECT 143.100 43.400 144.900 43.700 ;
        RECT 143.500 43.100 143.800 43.400 ;
        RECT 146.200 43.100 146.600 43.500 ;
        RECT 141.100 41.100 141.700 43.100 ;
        RECT 143.400 41.100 143.800 43.100 ;
        RECT 145.600 42.800 146.600 43.100 ;
        RECT 145.600 41.100 146.000 42.800 ;
        RECT 147.800 41.100 148.200 45.300 ;
        RECT 151.100 45.100 151.400 46.800 ;
        RECT 152.600 46.800 153.000 47.200 ;
        RECT 153.400 46.800 153.800 47.200 ;
        RECT 155.600 49.100 156.000 49.900 ;
        RECT 156.600 49.100 157.000 49.200 ;
        RECT 155.600 48.800 157.000 49.100 ;
        RECT 155.600 47.100 156.000 48.800 ;
        RECT 151.800 45.400 152.200 46.200 ;
        RECT 152.600 46.100 152.900 46.800 ;
        RECT 153.500 46.100 153.800 46.800 ;
        RECT 155.100 46.900 156.000 47.100 ;
        RECT 158.200 47.700 158.600 49.900 ;
        RECT 160.300 49.200 160.900 49.900 ;
        RECT 160.300 48.900 161.000 49.200 ;
        RECT 162.600 48.900 163.000 49.900 ;
        RECT 164.800 49.200 165.200 49.900 ;
        RECT 164.800 48.900 165.800 49.200 ;
        RECT 160.600 48.500 161.000 48.900 ;
        RECT 162.700 48.600 163.000 48.900 ;
        RECT 162.700 48.300 164.100 48.600 ;
        RECT 163.700 48.200 164.100 48.300 ;
        RECT 164.600 48.200 165.000 48.600 ;
        RECT 165.400 48.500 165.800 48.900 ;
        RECT 159.700 47.700 160.100 47.800 ;
        RECT 158.200 47.400 160.100 47.700 ;
        RECT 155.100 46.800 155.900 46.900 ;
        RECT 152.600 45.800 153.800 46.100 ;
        RECT 153.500 45.100 153.800 45.800 ;
        RECT 154.200 45.400 154.600 46.200 ;
        RECT 155.100 45.200 155.400 46.800 ;
        RECT 156.200 45.800 157.000 46.200 ;
        RECT 158.200 45.700 158.600 47.400 ;
        RECT 161.700 47.100 162.100 47.200 ;
        RECT 164.600 47.100 164.900 48.200 ;
        RECT 167.000 47.500 167.400 49.900 ;
        RECT 168.100 48.200 168.500 49.900 ;
        RECT 171.000 48.900 171.400 49.900 ;
        RECT 168.100 47.900 169.000 48.200 ;
        RECT 166.200 47.100 167.000 47.200 ;
        RECT 161.500 46.800 167.000 47.100 ;
        RECT 160.600 46.400 161.000 46.500 ;
        RECT 159.100 46.100 161.000 46.400 ;
        RECT 159.100 46.000 159.500 46.100 ;
        RECT 159.900 45.700 160.300 45.800 ;
        RECT 151.000 44.700 151.900 45.100 ;
        RECT 153.400 44.700 154.300 45.100 ;
        RECT 155.000 44.800 155.400 45.200 ;
        RECT 157.400 44.800 157.800 45.600 ;
        RECT 158.200 45.400 160.300 45.700 ;
        RECT 151.500 41.100 151.900 44.700 ;
        RECT 153.900 41.100 154.300 44.700 ;
        RECT 155.100 43.500 155.400 44.800 ;
        RECT 155.800 43.800 156.200 44.600 ;
        RECT 155.100 43.200 156.900 43.500 ;
        RECT 155.100 43.100 155.400 43.200 ;
        RECT 155.000 41.100 155.400 43.100 ;
        RECT 156.600 43.100 156.900 43.200 ;
        RECT 156.600 41.100 157.000 43.100 ;
        RECT 158.200 41.100 158.600 45.400 ;
        RECT 161.500 45.200 161.800 46.800 ;
        RECT 165.100 46.700 165.500 46.800 ;
        RECT 164.600 46.200 165.000 46.300 ;
        RECT 165.900 46.200 166.300 46.300 ;
        RECT 163.800 45.900 166.300 46.200 ;
        RECT 163.800 45.800 164.200 45.900 ;
        RECT 164.600 45.500 167.400 45.600 ;
        RECT 164.500 45.400 167.400 45.500 ;
        RECT 160.600 44.900 161.800 45.200 ;
        RECT 162.500 45.300 167.400 45.400 ;
        RECT 162.500 45.100 164.900 45.300 ;
        RECT 160.600 44.400 160.900 44.900 ;
        RECT 160.200 44.200 160.900 44.400 ;
        RECT 161.700 44.500 162.100 44.600 ;
        RECT 162.500 44.500 162.800 45.100 ;
        RECT 161.700 44.200 162.800 44.500 ;
        RECT 163.100 44.500 165.800 44.800 ;
        RECT 163.100 44.400 163.500 44.500 ;
        RECT 165.400 44.400 165.800 44.500 ;
        RECT 159.800 44.000 160.900 44.200 ;
        RECT 159.800 43.800 160.500 44.000 ;
        RECT 162.300 43.700 162.700 43.800 ;
        RECT 163.700 43.700 164.100 43.800 ;
        RECT 160.600 43.100 161.000 43.500 ;
        RECT 162.300 43.400 164.100 43.700 ;
        RECT 162.700 43.100 163.000 43.400 ;
        RECT 165.400 43.100 165.800 43.500 ;
        RECT 160.300 41.100 160.900 43.100 ;
        RECT 162.600 41.100 163.000 43.100 ;
        RECT 164.800 42.800 165.800 43.100 ;
        RECT 164.800 41.100 165.200 42.800 ;
        RECT 167.000 41.100 167.400 45.300 ;
        RECT 167.800 44.400 168.200 45.200 ;
        RECT 168.600 41.100 169.000 47.900 ;
        RECT 170.200 47.800 170.600 48.600 ;
        RECT 169.400 46.800 169.800 47.600 ;
        RECT 171.100 47.200 171.400 48.900 ;
        RECT 172.600 47.500 173.000 49.900 ;
        RECT 174.800 49.200 175.200 49.900 ;
        RECT 174.200 48.900 175.200 49.200 ;
        RECT 177.000 48.900 177.400 49.900 ;
        RECT 179.100 49.200 179.700 49.900 ;
        RECT 179.000 48.900 179.700 49.200 ;
        RECT 174.200 48.500 174.600 48.900 ;
        RECT 177.000 48.600 177.300 48.900 ;
        RECT 175.000 48.200 175.400 48.600 ;
        RECT 175.900 48.300 177.300 48.600 ;
        RECT 179.000 48.500 179.400 48.900 ;
        RECT 175.900 48.200 176.300 48.300 ;
        RECT 171.000 46.800 171.400 47.200 ;
        RECT 173.000 47.100 173.800 47.200 ;
        RECT 175.100 47.100 175.400 48.200 ;
        RECT 179.900 47.700 180.300 47.800 ;
        RECT 181.400 47.700 181.800 49.900 ;
        RECT 179.900 47.400 181.800 47.700 ;
        RECT 182.200 47.500 182.600 49.900 ;
        RECT 184.400 49.200 184.800 49.900 ;
        RECT 183.800 48.900 184.800 49.200 ;
        RECT 186.600 48.900 187.000 49.900 ;
        RECT 188.700 49.200 189.300 49.900 ;
        RECT 188.600 48.900 189.300 49.200 ;
        RECT 183.800 48.500 184.200 48.900 ;
        RECT 186.600 48.600 186.900 48.900 ;
        RECT 184.600 48.200 185.000 48.600 ;
        RECT 185.500 48.300 186.900 48.600 ;
        RECT 188.600 48.500 189.000 48.900 ;
        RECT 185.500 48.200 185.900 48.300 ;
        RECT 177.900 47.100 178.300 47.200 ;
        RECT 173.000 46.800 178.500 47.100 ;
        RECT 170.200 46.100 170.600 46.200 ;
        RECT 171.100 46.100 171.400 46.800 ;
        RECT 174.500 46.700 174.900 46.800 ;
        RECT 173.700 46.200 174.100 46.300 ;
        RECT 175.000 46.200 175.400 46.300 ;
        RECT 170.200 45.800 171.400 46.100 ;
        RECT 171.100 45.100 171.400 45.800 ;
        RECT 171.800 45.400 172.200 46.200 ;
        RECT 173.700 45.900 176.200 46.200 ;
        RECT 175.800 45.800 176.200 45.900 ;
        RECT 172.600 45.500 175.400 45.600 ;
        RECT 172.600 45.400 175.500 45.500 ;
        RECT 172.600 45.300 177.500 45.400 ;
        RECT 171.000 44.700 171.900 45.100 ;
        RECT 171.500 41.100 171.900 44.700 ;
        RECT 172.600 41.100 173.000 45.300 ;
        RECT 175.100 45.100 177.500 45.300 ;
        RECT 174.200 44.500 176.900 44.800 ;
        RECT 174.200 44.400 174.600 44.500 ;
        RECT 176.500 44.400 176.900 44.500 ;
        RECT 177.200 44.500 177.500 45.100 ;
        RECT 178.200 45.200 178.500 46.800 ;
        RECT 179.000 46.400 179.400 46.500 ;
        RECT 179.000 46.100 180.900 46.400 ;
        RECT 180.500 46.000 180.900 46.100 ;
        RECT 179.700 45.700 180.100 45.800 ;
        RECT 181.400 45.700 181.800 47.400 ;
        RECT 182.600 47.100 183.400 47.200 ;
        RECT 184.700 47.100 185.000 48.200 ;
        RECT 189.500 47.700 189.900 47.800 ;
        RECT 191.000 47.700 191.400 49.900 ;
        RECT 189.500 47.400 191.400 47.700 ;
        RECT 187.500 47.100 187.900 47.200 ;
        RECT 182.600 46.800 188.100 47.100 ;
        RECT 184.100 46.700 184.500 46.800 ;
        RECT 183.300 46.200 183.700 46.300 ;
        RECT 183.300 45.900 185.800 46.200 ;
        RECT 185.400 45.800 185.800 45.900 ;
        RECT 187.000 46.100 187.400 46.200 ;
        RECT 187.800 46.100 188.100 46.800 ;
        RECT 188.600 46.400 189.000 46.500 ;
        RECT 188.600 46.100 190.500 46.400 ;
        RECT 187.000 45.800 188.100 46.100 ;
        RECT 190.100 46.000 190.500 46.100 ;
        RECT 179.700 45.400 181.800 45.700 ;
        RECT 178.200 44.900 179.400 45.200 ;
        RECT 177.900 44.500 178.300 44.600 ;
        RECT 177.200 44.200 178.300 44.500 ;
        RECT 179.100 44.400 179.400 44.900 ;
        RECT 179.100 44.000 179.800 44.400 ;
        RECT 175.900 43.700 176.300 43.800 ;
        RECT 177.300 43.700 177.700 43.800 ;
        RECT 174.200 43.100 174.600 43.500 ;
        RECT 175.900 43.400 177.700 43.700 ;
        RECT 177.000 43.100 177.300 43.400 ;
        RECT 179.000 43.100 179.400 43.500 ;
        RECT 174.200 42.800 175.200 43.100 ;
        RECT 174.800 41.100 175.200 42.800 ;
        RECT 177.000 41.100 177.400 43.100 ;
        RECT 179.100 41.100 179.700 43.100 ;
        RECT 181.400 41.100 181.800 45.400 ;
        RECT 182.200 45.500 185.000 45.600 ;
        RECT 182.200 45.400 185.100 45.500 ;
        RECT 182.200 45.300 187.100 45.400 ;
        RECT 182.200 41.100 182.600 45.300 ;
        RECT 184.700 45.100 187.100 45.300 ;
        RECT 183.800 44.500 186.500 44.800 ;
        RECT 183.800 44.400 184.200 44.500 ;
        RECT 186.100 44.400 186.500 44.500 ;
        RECT 186.800 44.500 187.100 45.100 ;
        RECT 187.800 45.200 188.100 45.800 ;
        RECT 189.300 45.700 189.700 45.800 ;
        RECT 191.000 45.700 191.400 47.400 ;
        RECT 191.800 47.600 192.200 49.900 ;
        RECT 191.800 47.300 192.900 47.600 ;
        RECT 189.300 45.400 191.400 45.700 ;
        RECT 187.800 44.900 189.000 45.200 ;
        RECT 187.500 44.500 187.900 44.600 ;
        RECT 186.800 44.200 187.900 44.500 ;
        RECT 188.700 44.400 189.000 44.900 ;
        RECT 188.700 44.000 189.400 44.400 ;
        RECT 185.500 43.700 185.900 43.800 ;
        RECT 186.900 43.700 187.300 43.800 ;
        RECT 183.800 43.100 184.200 43.500 ;
        RECT 185.500 43.400 187.300 43.700 ;
        RECT 186.600 43.100 186.900 43.400 ;
        RECT 188.600 43.100 189.000 43.500 ;
        RECT 183.800 42.800 184.800 43.100 ;
        RECT 184.400 41.100 184.800 42.800 ;
        RECT 186.600 41.100 187.000 43.100 ;
        RECT 188.700 41.100 189.300 43.100 ;
        RECT 191.000 41.100 191.400 45.400 ;
        RECT 192.600 45.800 192.900 47.300 ;
        RECT 193.400 46.200 193.800 49.900 ;
        RECT 192.600 45.400 193.200 45.800 ;
        RECT 192.600 45.100 192.900 45.400 ;
        RECT 193.500 45.100 193.800 46.200 ;
        RECT 191.800 44.800 192.900 45.100 ;
        RECT 191.800 41.100 192.200 44.800 ;
        RECT 193.400 41.100 193.800 45.100 ;
        RECT 0.600 35.600 1.000 39.900 ;
        RECT 2.700 37.900 3.300 39.900 ;
        RECT 5.000 37.900 5.400 39.900 ;
        RECT 7.200 38.200 7.600 39.900 ;
        RECT 7.200 37.900 8.200 38.200 ;
        RECT 3.000 37.500 3.400 37.900 ;
        RECT 5.100 37.600 5.400 37.900 ;
        RECT 4.700 37.300 6.500 37.600 ;
        RECT 7.800 37.500 8.200 37.900 ;
        RECT 4.700 37.200 5.100 37.300 ;
        RECT 6.100 37.200 6.500 37.300 ;
        RECT 2.600 36.600 3.300 37.000 ;
        RECT 3.000 36.100 3.300 36.600 ;
        RECT 4.100 36.500 5.200 36.800 ;
        RECT 4.100 36.400 4.500 36.500 ;
        RECT 3.000 35.800 4.200 36.100 ;
        RECT 0.600 35.300 2.700 35.600 ;
        RECT 0.600 33.600 1.000 35.300 ;
        RECT 2.300 35.200 2.700 35.300 ;
        RECT 1.500 34.900 1.900 35.000 ;
        RECT 1.500 34.600 3.400 34.900 ;
        RECT 3.000 34.500 3.400 34.600 ;
        RECT 3.900 34.200 4.200 35.800 ;
        RECT 4.900 35.900 5.200 36.500 ;
        RECT 5.500 36.500 5.900 36.600 ;
        RECT 7.800 36.500 8.200 36.600 ;
        RECT 5.500 36.200 8.200 36.500 ;
        RECT 4.900 35.700 7.300 35.900 ;
        RECT 9.400 35.700 9.800 39.900 ;
        RECT 4.900 35.600 9.800 35.700 ;
        RECT 6.900 35.500 9.800 35.600 ;
        RECT 7.000 35.400 9.800 35.500 ;
        RECT 10.200 35.600 10.600 39.900 ;
        RECT 12.300 37.900 12.900 39.900 ;
        RECT 14.600 37.900 15.000 39.900 ;
        RECT 16.800 38.200 17.200 39.900 ;
        RECT 16.800 37.900 17.800 38.200 ;
        RECT 12.600 37.500 13.000 37.900 ;
        RECT 14.700 37.600 15.000 37.900 ;
        RECT 14.300 37.300 16.100 37.600 ;
        RECT 17.400 37.500 17.800 37.900 ;
        RECT 14.300 37.200 14.700 37.300 ;
        RECT 15.700 37.200 16.100 37.300 ;
        RECT 12.200 36.600 12.900 37.000 ;
        RECT 12.600 36.100 12.900 36.600 ;
        RECT 13.700 36.500 14.800 36.800 ;
        RECT 13.700 36.400 14.100 36.500 ;
        RECT 12.600 35.800 13.800 36.100 ;
        RECT 10.200 35.300 12.300 35.600 ;
        RECT 6.200 35.100 6.600 35.200 ;
        RECT 6.200 34.800 8.700 35.100 ;
        RECT 7.000 34.700 7.400 34.800 ;
        RECT 8.300 34.700 8.700 34.800 ;
        RECT 7.500 34.200 7.900 34.300 ;
        RECT 3.900 33.900 9.400 34.200 ;
        RECT 4.100 33.800 4.500 33.900 ;
        RECT 0.600 33.300 2.500 33.600 ;
        RECT 0.600 31.100 1.000 33.300 ;
        RECT 2.100 33.200 2.500 33.300 ;
        RECT 7.000 32.800 7.300 33.900 ;
        RECT 8.600 33.800 9.400 33.900 ;
        RECT 10.200 33.600 10.600 35.300 ;
        RECT 11.900 35.200 12.300 35.300 ;
        RECT 11.100 34.900 11.500 35.000 ;
        RECT 11.100 34.600 13.000 34.900 ;
        RECT 12.600 34.500 13.000 34.600 ;
        RECT 13.500 34.200 13.800 35.800 ;
        RECT 14.500 35.900 14.800 36.500 ;
        RECT 15.100 36.500 15.500 36.600 ;
        RECT 17.400 36.500 17.800 36.600 ;
        RECT 15.100 36.200 17.800 36.500 ;
        RECT 14.500 35.700 16.900 35.900 ;
        RECT 19.000 35.700 19.400 39.900 ;
        RECT 14.500 35.600 19.400 35.700 ;
        RECT 16.500 35.500 19.400 35.600 ;
        RECT 16.600 35.400 19.400 35.500 ;
        RECT 19.800 35.700 20.200 39.900 ;
        RECT 22.000 38.200 22.400 39.900 ;
        RECT 21.400 37.900 22.400 38.200 ;
        RECT 24.200 37.900 24.600 39.900 ;
        RECT 26.300 37.900 26.900 39.900 ;
        RECT 21.400 37.500 21.800 37.900 ;
        RECT 24.200 37.600 24.500 37.900 ;
        RECT 23.100 37.300 24.900 37.600 ;
        RECT 26.200 37.500 26.600 37.900 ;
        RECT 23.100 37.200 23.500 37.300 ;
        RECT 24.500 37.200 24.900 37.300 ;
        RECT 21.400 36.500 21.800 36.600 ;
        RECT 23.700 36.500 24.100 36.600 ;
        RECT 21.400 36.200 24.100 36.500 ;
        RECT 24.400 36.500 25.500 36.800 ;
        RECT 24.400 35.900 24.700 36.500 ;
        RECT 25.100 36.400 25.500 36.500 ;
        RECT 26.300 36.600 27.000 37.000 ;
        RECT 26.300 36.100 26.600 36.600 ;
        RECT 22.300 35.700 24.700 35.900 ;
        RECT 19.800 35.600 24.700 35.700 ;
        RECT 25.400 35.800 26.600 36.100 ;
        RECT 19.800 35.500 22.700 35.600 ;
        RECT 19.800 35.400 22.600 35.500 ;
        RECT 14.200 35.100 14.600 35.200 ;
        RECT 15.800 35.100 16.200 35.200 ;
        RECT 23.000 35.100 23.400 35.200 ;
        RECT 14.200 34.800 18.300 35.100 ;
        RECT 17.900 34.700 18.300 34.800 ;
        RECT 20.900 34.800 23.400 35.100 ;
        RECT 20.900 34.700 21.300 34.800 ;
        RECT 22.200 34.700 22.600 34.800 ;
        RECT 17.100 34.200 17.500 34.300 ;
        RECT 21.700 34.200 22.100 34.300 ;
        RECT 25.400 34.200 25.700 35.800 ;
        RECT 28.600 35.600 29.000 39.900 ;
        RECT 26.900 35.300 29.000 35.600 ;
        RECT 26.900 35.200 27.300 35.300 ;
        RECT 27.700 34.900 28.100 35.000 ;
        RECT 26.200 34.600 28.100 34.900 ;
        RECT 26.200 34.500 26.600 34.600 ;
        RECT 13.500 34.100 19.000 34.200 ;
        RECT 20.200 34.100 25.700 34.200 ;
        RECT 13.500 33.900 25.700 34.100 ;
        RECT 13.700 33.800 14.100 33.900 ;
        RECT 6.100 32.700 6.500 32.800 ;
        RECT 3.000 32.100 3.400 32.500 ;
        RECT 5.100 32.400 6.500 32.700 ;
        RECT 7.000 32.400 7.400 32.800 ;
        RECT 5.100 32.100 5.400 32.400 ;
        RECT 7.800 32.100 8.200 32.500 ;
        RECT 2.700 31.800 3.400 32.100 ;
        RECT 2.700 31.100 3.300 31.800 ;
        RECT 5.000 31.100 5.400 32.100 ;
        RECT 7.200 31.800 8.200 32.100 ;
        RECT 7.200 31.100 7.600 31.800 ;
        RECT 9.400 31.100 9.800 33.500 ;
        RECT 10.200 33.300 12.100 33.600 ;
        RECT 10.200 31.100 10.600 33.300 ;
        RECT 11.700 33.200 12.100 33.300 ;
        RECT 16.600 32.800 16.900 33.900 ;
        RECT 18.200 33.800 21.000 33.900 ;
        RECT 15.700 32.700 16.100 32.800 ;
        RECT 12.600 32.100 13.000 32.500 ;
        RECT 14.700 32.400 16.100 32.700 ;
        RECT 16.600 32.400 17.000 32.800 ;
        RECT 14.700 32.100 15.000 32.400 ;
        RECT 17.400 32.100 17.800 32.500 ;
        RECT 12.300 31.800 13.000 32.100 ;
        RECT 12.300 31.100 12.900 31.800 ;
        RECT 14.600 31.100 15.000 32.100 ;
        RECT 16.800 31.800 17.800 32.100 ;
        RECT 16.800 31.100 17.200 31.800 ;
        RECT 19.000 31.100 19.400 33.500 ;
        RECT 19.800 31.100 20.200 33.500 ;
        RECT 22.300 32.800 22.600 33.900 ;
        RECT 23.800 33.800 24.200 33.900 ;
        RECT 25.100 33.800 25.500 33.900 ;
        RECT 28.600 33.600 29.000 35.300 ;
        RECT 27.100 33.300 29.000 33.600 ;
        RECT 27.100 33.200 27.500 33.300 ;
        RECT 21.400 32.100 21.800 32.500 ;
        RECT 22.200 32.400 22.600 32.800 ;
        RECT 23.100 32.700 23.500 32.800 ;
        RECT 23.100 32.400 24.500 32.700 ;
        RECT 24.200 32.100 24.500 32.400 ;
        RECT 26.200 32.100 26.600 32.500 ;
        RECT 21.400 31.800 22.400 32.100 ;
        RECT 22.000 31.100 22.400 31.800 ;
        RECT 24.200 31.100 24.600 32.100 ;
        RECT 26.200 31.800 26.900 32.100 ;
        RECT 26.300 31.100 26.900 31.800 ;
        RECT 28.600 31.100 29.000 33.300 ;
        RECT 29.400 35.600 29.800 39.900 ;
        RECT 31.500 37.900 32.100 39.900 ;
        RECT 33.800 37.900 34.200 39.900 ;
        RECT 36.000 38.200 36.400 39.900 ;
        RECT 36.000 37.900 37.000 38.200 ;
        RECT 31.800 37.500 32.200 37.900 ;
        RECT 33.900 37.600 34.200 37.900 ;
        RECT 33.500 37.300 35.300 37.600 ;
        RECT 36.600 37.500 37.000 37.900 ;
        RECT 33.500 37.200 33.900 37.300 ;
        RECT 34.900 37.200 35.300 37.300 ;
        RECT 31.400 36.600 32.100 37.000 ;
        RECT 31.800 36.100 32.100 36.600 ;
        RECT 32.900 36.500 34.000 36.800 ;
        RECT 32.900 36.400 33.300 36.500 ;
        RECT 31.800 35.800 33.000 36.100 ;
        RECT 29.400 35.300 31.500 35.600 ;
        RECT 29.400 33.600 29.800 35.300 ;
        RECT 31.100 35.200 31.500 35.300 ;
        RECT 30.300 34.900 30.700 35.000 ;
        RECT 30.300 34.600 32.200 34.900 ;
        RECT 31.800 34.500 32.200 34.600 ;
        RECT 32.700 34.200 33.000 35.800 ;
        RECT 33.700 35.900 34.000 36.500 ;
        RECT 34.300 36.500 34.700 36.600 ;
        RECT 36.600 36.500 37.000 36.600 ;
        RECT 34.300 36.200 37.000 36.500 ;
        RECT 33.700 35.700 36.100 35.900 ;
        RECT 38.200 35.700 38.600 39.900 ;
        RECT 39.800 37.900 40.200 39.900 ;
        RECT 33.700 35.600 38.600 35.700 ;
        RECT 35.700 35.500 38.600 35.600 ;
        RECT 39.900 35.800 40.200 37.900 ;
        RECT 41.400 35.900 41.800 39.900 ;
        RECT 43.500 39.200 44.500 39.900 ;
        RECT 43.000 38.800 44.500 39.200 ;
        RECT 43.500 35.900 44.500 38.800 ;
        RECT 47.800 35.900 48.200 39.900 ;
        RECT 49.400 37.900 49.800 39.900 ;
        RECT 39.900 35.500 41.100 35.800 ;
        RECT 35.800 35.400 38.600 35.500 ;
        RECT 35.000 35.100 35.400 35.200 ;
        RECT 35.000 34.800 37.500 35.100 ;
        RECT 39.800 34.800 40.200 35.200 ;
        RECT 35.800 34.700 36.200 34.800 ;
        RECT 37.100 34.700 37.500 34.800 ;
        RECT 36.300 34.200 36.700 34.300 ;
        RECT 32.600 33.900 38.200 34.200 ;
        RECT 32.600 33.800 33.300 33.900 ;
        RECT 29.400 33.300 31.300 33.600 ;
        RECT 29.400 31.100 29.800 33.300 ;
        RECT 30.900 33.200 31.300 33.300 ;
        RECT 32.600 33.200 32.900 33.800 ;
        RECT 35.800 33.200 36.100 33.900 ;
        RECT 37.400 33.800 38.200 33.900 ;
        RECT 39.000 33.800 39.400 34.600 ;
        RECT 39.900 34.400 40.200 34.800 ;
        RECT 39.900 34.100 40.400 34.400 ;
        RECT 40.000 34.000 40.400 34.100 ;
        RECT 40.800 33.800 41.100 35.500 ;
        RECT 41.500 35.200 41.800 35.900 ;
        RECT 41.400 35.100 41.800 35.200 ;
        RECT 41.400 34.800 42.500 35.100 ;
        RECT 40.800 33.700 41.200 33.800 ;
        RECT 39.700 33.500 41.200 33.700 ;
        RECT 32.600 32.800 33.000 33.200 ;
        RECT 34.900 32.700 35.300 32.800 ;
        RECT 31.800 32.100 32.200 32.500 ;
        RECT 33.900 32.400 35.300 32.700 ;
        RECT 35.800 32.400 36.200 33.200 ;
        RECT 33.900 32.100 34.200 32.400 ;
        RECT 36.600 32.100 37.000 32.500 ;
        RECT 31.500 31.800 32.200 32.100 ;
        RECT 31.500 31.100 32.100 31.800 ;
        RECT 33.800 31.100 34.200 32.100 ;
        RECT 36.000 31.800 37.000 32.100 ;
        RECT 36.000 31.100 36.400 31.800 ;
        RECT 38.200 31.100 38.600 33.500 ;
        RECT 39.100 33.400 41.200 33.500 ;
        RECT 39.100 33.200 40.000 33.400 ;
        RECT 39.100 33.100 39.400 33.200 ;
        RECT 41.500 33.100 41.800 34.800 ;
        RECT 42.200 34.200 42.500 34.800 ;
        RECT 43.000 34.400 43.400 35.200 ;
        RECT 43.800 34.200 44.100 35.900 ;
        RECT 47.800 35.200 48.100 35.900 ;
        RECT 49.400 35.800 49.700 37.900 ;
        RECT 51.300 36.300 51.700 39.900 ;
        RECT 51.300 35.900 52.200 36.300 ;
        RECT 48.500 35.500 49.700 35.800 ;
        RECT 44.600 34.400 45.000 35.200 ;
        RECT 47.800 35.100 48.200 35.200 ;
        RECT 46.200 34.800 48.200 35.100 ;
        RECT 42.200 34.100 42.600 34.200 ;
        RECT 43.800 34.100 44.200 34.200 ;
        RECT 45.400 34.100 45.800 34.600 ;
        RECT 46.200 34.100 46.500 34.800 ;
        RECT 42.200 33.800 43.000 34.100 ;
        RECT 43.800 33.800 45.000 34.100 ;
        RECT 45.400 33.800 46.500 34.100 ;
        RECT 42.600 33.600 43.000 33.800 ;
        RECT 42.300 33.100 44.100 33.300 ;
        RECT 44.700 33.100 45.000 33.800 ;
        RECT 47.800 33.100 48.100 34.800 ;
        RECT 48.500 33.800 48.800 35.500 ;
        RECT 49.400 34.800 49.800 35.200 ;
        RECT 51.000 34.800 51.400 35.600 ;
        RECT 51.800 35.100 52.100 35.900 ;
        RECT 53.400 35.600 53.800 39.900 ;
        RECT 55.500 37.900 56.100 39.900 ;
        RECT 57.800 37.900 58.200 39.900 ;
        RECT 60.000 38.200 60.400 39.900 ;
        RECT 60.000 37.900 61.000 38.200 ;
        RECT 55.800 37.500 56.200 37.900 ;
        RECT 57.900 37.600 58.200 37.900 ;
        RECT 57.500 37.300 59.300 37.600 ;
        RECT 60.600 37.500 61.000 37.900 ;
        RECT 57.500 37.200 57.900 37.300 ;
        RECT 58.900 37.200 59.300 37.300 ;
        RECT 55.400 36.600 56.100 37.000 ;
        RECT 55.800 36.100 56.100 36.600 ;
        RECT 56.900 36.500 58.000 36.800 ;
        RECT 56.900 36.400 57.300 36.500 ;
        RECT 55.800 35.800 57.000 36.100 ;
        RECT 53.400 35.300 55.500 35.600 ;
        RECT 52.600 35.100 53.000 35.200 ;
        RECT 51.800 34.800 53.000 35.100 ;
        RECT 49.400 34.400 49.700 34.800 ;
        RECT 49.200 34.100 49.700 34.400 ;
        RECT 49.200 34.000 49.600 34.100 ;
        RECT 50.200 33.800 50.600 34.600 ;
        RECT 51.800 34.200 52.100 34.800 ;
        RECT 51.800 33.800 52.200 34.200 ;
        RECT 48.400 33.700 48.800 33.800 ;
        RECT 48.400 33.500 49.900 33.700 ;
        RECT 48.400 33.400 50.500 33.500 ;
        RECT 49.600 33.200 50.500 33.400 ;
        RECT 50.200 33.100 50.500 33.200 ;
        RECT 39.000 31.100 39.400 33.100 ;
        RECT 41.100 32.600 41.800 33.100 ;
        RECT 42.200 33.000 44.200 33.100 ;
        RECT 41.100 31.100 41.500 32.600 ;
        RECT 42.200 31.100 42.600 33.000 ;
        RECT 43.800 31.400 44.200 33.000 ;
        RECT 44.600 31.700 45.000 33.100 ;
        RECT 45.400 31.400 45.800 33.100 ;
        RECT 47.800 32.600 48.500 33.100 ;
        RECT 43.800 31.100 45.800 31.400 ;
        RECT 48.100 31.100 48.500 32.600 ;
        RECT 50.200 31.100 50.600 33.100 ;
        RECT 51.800 32.100 52.100 33.800 ;
        RECT 53.400 33.600 53.800 35.300 ;
        RECT 55.100 35.200 55.500 35.300 ;
        RECT 56.700 35.100 57.000 35.800 ;
        RECT 57.700 35.900 58.000 36.500 ;
        RECT 58.300 36.500 58.700 36.600 ;
        RECT 60.600 36.500 61.000 36.600 ;
        RECT 58.300 36.200 61.000 36.500 ;
        RECT 57.700 35.700 60.100 35.900 ;
        RECT 62.200 35.700 62.600 39.900 ;
        RECT 63.300 36.200 63.700 39.900 ;
        RECT 57.700 35.600 62.600 35.700 ;
        RECT 59.700 35.500 62.600 35.600 ;
        RECT 59.800 35.400 62.600 35.500 ;
        RECT 63.000 35.900 63.700 36.200 ;
        RECT 63.000 35.200 63.300 35.900 ;
        RECT 65.400 35.600 65.800 39.900 ;
        RECT 63.800 35.400 65.800 35.600 ;
        RECT 63.700 35.300 65.800 35.400 ;
        RECT 57.400 35.100 57.800 35.200 ;
        RECT 54.300 34.900 54.700 35.000 ;
        RECT 54.300 34.600 56.200 34.900 ;
        RECT 56.600 34.800 57.800 35.100 ;
        RECT 59.000 35.100 59.400 35.200 ;
        RECT 59.000 34.800 61.500 35.100 ;
        RECT 55.800 34.500 56.200 34.600 ;
        RECT 56.700 34.200 57.000 34.800 ;
        RECT 59.800 34.700 60.200 34.800 ;
        RECT 61.100 34.700 61.500 34.800 ;
        RECT 63.000 34.800 63.400 35.200 ;
        RECT 63.700 35.000 64.100 35.300 ;
        RECT 67.000 35.100 67.400 39.900 ;
        RECT 69.100 36.300 69.500 39.900 ;
        RECT 68.600 35.900 69.500 36.300 ;
        RECT 60.300 34.200 60.700 34.300 ;
        RECT 54.200 33.600 54.600 34.200 ;
        RECT 56.700 33.900 62.200 34.200 ;
        RECT 56.900 33.800 57.300 33.900 ;
        RECT 53.400 33.300 55.300 33.600 ;
        RECT 52.600 32.400 53.000 33.200 ;
        RECT 51.800 31.100 52.200 32.100 ;
        RECT 53.400 31.100 53.800 33.300 ;
        RECT 54.900 33.200 55.300 33.300 ;
        RECT 59.800 32.800 60.100 33.900 ;
        RECT 61.400 33.800 62.200 33.900 ;
        RECT 58.900 32.700 59.300 32.800 ;
        RECT 55.800 32.100 56.200 32.500 ;
        RECT 57.900 32.400 59.300 32.700 ;
        RECT 59.800 32.400 60.200 32.800 ;
        RECT 57.900 32.100 58.200 32.400 ;
        RECT 60.600 32.100 61.000 32.500 ;
        RECT 55.500 31.800 56.200 32.100 ;
        RECT 55.500 31.100 56.100 31.800 ;
        RECT 57.800 31.100 58.200 32.100 ;
        RECT 60.000 31.800 61.000 32.100 ;
        RECT 60.000 31.100 60.400 31.800 ;
        RECT 62.200 31.100 62.600 33.500 ;
        RECT 63.000 33.100 63.300 34.800 ;
        RECT 63.700 33.500 64.000 35.000 ;
        RECT 67.000 34.800 68.100 35.100 ;
        RECT 64.400 34.200 64.800 34.600 ;
        RECT 64.500 33.800 65.000 34.200 ;
        RECT 63.700 33.200 64.900 33.500 ;
        RECT 63.000 31.100 63.400 33.100 ;
        RECT 64.600 32.100 64.900 33.200 ;
        RECT 66.200 32.400 66.600 33.200 ;
        RECT 64.600 31.100 65.000 32.100 ;
        RECT 67.000 31.100 67.400 34.800 ;
        RECT 67.800 34.200 68.100 34.800 ;
        RECT 68.700 34.200 69.000 35.900 ;
        RECT 70.200 35.800 70.600 36.600 ;
        RECT 69.400 35.100 69.800 35.600 ;
        RECT 70.200 35.100 70.500 35.800 ;
        RECT 69.400 34.800 70.500 35.100 ;
        RECT 67.800 33.800 68.200 34.200 ;
        RECT 68.600 33.800 69.000 34.200 ;
        RECT 68.700 32.100 69.000 33.800 ;
        RECT 71.000 33.100 71.400 39.900 ;
        RECT 72.600 35.900 73.000 39.900 ;
        RECT 74.200 37.900 74.600 39.900 ;
        RECT 72.600 35.200 72.900 35.900 ;
        RECT 74.200 35.800 74.500 37.900 ;
        RECT 77.100 36.300 77.500 39.900 ;
        RECT 78.200 37.100 78.600 37.200 ;
        RECT 79.000 37.100 79.400 39.900 ;
        RECT 78.200 36.800 79.400 37.100 ;
        RECT 76.600 35.900 77.500 36.300 ;
        RECT 73.300 35.500 74.500 35.800 ;
        RECT 72.600 34.800 73.000 35.200 ;
        RECT 71.800 33.400 72.200 34.200 ;
        RECT 68.600 31.100 69.000 32.100 ;
        RECT 70.500 32.800 71.400 33.100 ;
        RECT 72.600 33.100 72.900 34.800 ;
        RECT 73.300 33.800 73.600 35.500 ;
        RECT 74.200 34.800 74.600 35.200 ;
        RECT 74.200 34.400 74.500 34.800 ;
        RECT 74.000 34.100 74.500 34.400 ;
        RECT 74.000 34.000 74.400 34.100 ;
        RECT 75.000 33.800 75.400 34.600 ;
        RECT 76.700 34.200 77.000 35.900 ;
        RECT 77.400 35.100 77.800 35.600 ;
        RECT 79.000 35.100 79.400 36.800 ;
        RECT 79.800 35.700 80.200 39.900 ;
        RECT 82.000 38.200 82.400 39.900 ;
        RECT 81.400 37.900 82.400 38.200 ;
        RECT 84.200 37.900 84.600 39.900 ;
        RECT 86.300 37.900 86.900 39.900 ;
        RECT 81.400 37.500 81.800 37.900 ;
        RECT 84.200 37.600 84.500 37.900 ;
        RECT 83.100 37.300 84.900 37.600 ;
        RECT 86.200 37.500 86.600 37.900 ;
        RECT 83.100 37.200 83.500 37.300 ;
        RECT 84.500 37.200 84.900 37.300 ;
        RECT 81.400 36.500 81.800 36.600 ;
        RECT 83.700 36.500 84.100 36.600 ;
        RECT 81.400 36.200 84.100 36.500 ;
        RECT 84.400 36.500 85.500 36.800 ;
        RECT 84.400 35.900 84.700 36.500 ;
        RECT 85.100 36.400 85.500 36.500 ;
        RECT 86.300 36.600 87.000 37.000 ;
        RECT 86.300 36.100 86.600 36.600 ;
        RECT 82.300 35.700 84.700 35.900 ;
        RECT 79.800 35.600 84.700 35.700 ;
        RECT 85.400 35.800 86.600 36.100 ;
        RECT 79.800 35.500 82.700 35.600 ;
        RECT 79.800 35.400 82.600 35.500 ;
        RECT 83.000 35.100 83.400 35.200 ;
        RECT 84.600 35.100 85.000 35.200 ;
        RECT 77.400 34.800 79.400 35.100 ;
        RECT 76.600 33.800 77.000 34.200 ;
        RECT 73.200 33.700 73.600 33.800 ;
        RECT 73.200 33.500 74.700 33.700 ;
        RECT 73.200 33.400 75.300 33.500 ;
        RECT 74.400 33.200 75.300 33.400 ;
        RECT 75.000 33.100 75.300 33.200 ;
        RECT 70.500 31.100 70.900 32.800 ;
        RECT 72.600 32.600 73.300 33.100 ;
        RECT 72.900 31.100 73.300 32.600 ;
        RECT 75.000 31.100 75.400 33.100 ;
        RECT 76.700 32.100 77.000 33.800 ;
        RECT 78.200 32.400 78.600 33.200 ;
        RECT 76.600 31.100 77.000 32.100 ;
        RECT 79.000 31.100 79.400 34.800 ;
        RECT 80.900 34.800 85.000 35.100 ;
        RECT 80.900 34.700 81.300 34.800 ;
        RECT 81.700 34.200 82.100 34.300 ;
        RECT 85.400 34.200 85.700 35.800 ;
        RECT 88.600 35.600 89.000 39.900 ;
        RECT 86.900 35.300 89.000 35.600 ;
        RECT 89.400 35.700 89.800 39.900 ;
        RECT 91.600 38.200 92.000 39.900 ;
        RECT 91.000 37.900 92.000 38.200 ;
        RECT 93.800 37.900 94.200 39.900 ;
        RECT 95.900 37.900 96.500 39.900 ;
        RECT 98.200 39.100 98.600 39.900 ;
        RECT 99.800 39.100 100.200 39.200 ;
        RECT 98.200 38.800 100.200 39.100 ;
        RECT 91.000 37.500 91.400 37.900 ;
        RECT 93.800 37.600 94.100 37.900 ;
        RECT 92.700 37.300 94.500 37.600 ;
        RECT 95.800 37.500 96.200 37.900 ;
        RECT 92.700 37.200 93.100 37.300 ;
        RECT 94.100 37.200 94.500 37.300 ;
        RECT 91.000 36.500 91.400 36.600 ;
        RECT 93.300 36.500 93.700 36.600 ;
        RECT 91.000 36.200 93.700 36.500 ;
        RECT 94.000 36.500 95.100 36.800 ;
        RECT 94.000 35.900 94.300 36.500 ;
        RECT 94.700 36.400 95.100 36.500 ;
        RECT 95.900 36.600 96.600 37.000 ;
        RECT 95.900 36.100 96.200 36.600 ;
        RECT 91.900 35.700 94.300 35.900 ;
        RECT 89.400 35.600 94.300 35.700 ;
        RECT 95.000 35.800 96.200 36.100 ;
        RECT 89.400 35.500 92.300 35.600 ;
        RECT 89.400 35.400 92.200 35.500 ;
        RECT 86.900 35.200 87.300 35.300 ;
        RECT 87.700 34.900 88.100 35.000 ;
        RECT 86.200 34.600 88.100 34.900 ;
        RECT 86.200 34.500 86.600 34.600 ;
        RECT 80.200 33.900 85.700 34.200 ;
        RECT 80.200 33.800 81.000 33.900 ;
        RECT 79.800 31.100 80.200 33.500 ;
        RECT 82.300 32.800 82.600 33.900 ;
        RECT 83.800 33.800 84.200 33.900 ;
        RECT 85.100 33.800 85.500 33.900 ;
        RECT 88.600 33.600 89.000 35.300 ;
        RECT 92.600 35.100 93.000 35.200 ;
        RECT 90.500 34.800 93.000 35.100 ;
        RECT 90.500 34.700 90.900 34.800 ;
        RECT 91.800 34.700 92.200 34.800 ;
        RECT 91.300 34.200 91.700 34.300 ;
        RECT 95.000 34.200 95.300 35.800 ;
        RECT 98.200 35.600 98.600 38.800 ;
        RECT 96.500 35.300 98.600 35.600 ;
        RECT 96.500 35.200 96.900 35.300 ;
        RECT 97.300 34.900 97.700 35.000 ;
        RECT 95.800 34.600 97.700 34.900 ;
        RECT 95.800 34.500 96.200 34.600 ;
        RECT 89.800 33.900 95.300 34.200 ;
        RECT 89.800 33.800 90.600 33.900 ;
        RECT 87.100 33.300 89.000 33.600 ;
        RECT 87.100 33.200 87.500 33.300 ;
        RECT 81.400 32.100 81.800 32.500 ;
        RECT 82.200 32.400 82.600 32.800 ;
        RECT 83.100 32.700 83.500 32.800 ;
        RECT 83.100 32.400 84.500 32.700 ;
        RECT 84.200 32.100 84.500 32.400 ;
        RECT 86.200 32.100 86.600 32.500 ;
        RECT 81.400 31.800 82.400 32.100 ;
        RECT 82.000 31.100 82.400 31.800 ;
        RECT 84.200 31.100 84.600 32.100 ;
        RECT 86.200 31.800 86.900 32.100 ;
        RECT 86.300 31.100 86.900 31.800 ;
        RECT 88.600 31.100 89.000 33.300 ;
        RECT 89.400 31.100 89.800 33.500 ;
        RECT 91.900 33.200 92.200 33.900 ;
        RECT 94.700 33.800 95.100 33.900 ;
        RECT 98.200 33.600 98.600 35.300 ;
        RECT 96.700 33.300 98.600 33.600 ;
        RECT 96.700 33.200 97.100 33.300 ;
        RECT 91.000 32.100 91.400 32.500 ;
        RECT 91.800 32.400 92.200 33.200 ;
        RECT 92.700 32.700 93.100 32.800 ;
        RECT 92.700 32.400 94.100 32.700 ;
        RECT 93.800 32.100 94.100 32.400 ;
        RECT 95.800 32.100 96.200 32.500 ;
        RECT 91.000 31.800 92.000 32.100 ;
        RECT 91.600 31.100 92.000 31.800 ;
        RECT 93.800 31.100 94.200 32.100 ;
        RECT 95.800 31.800 96.500 32.100 ;
        RECT 95.900 31.100 96.500 31.800 ;
        RECT 98.200 31.100 98.600 33.300 ;
        RECT 100.600 35.900 101.000 39.900 ;
        RECT 102.200 37.900 102.600 39.900 ;
        RECT 100.600 35.200 100.900 35.900 ;
        RECT 102.200 35.800 102.500 37.900 ;
        RECT 103.800 36.900 104.200 39.900 ;
        RECT 103.900 36.600 104.200 36.900 ;
        RECT 105.400 39.600 107.400 39.900 ;
        RECT 105.400 36.900 105.800 39.600 ;
        RECT 106.200 36.900 106.600 39.300 ;
        RECT 107.000 37.000 107.400 39.600 ;
        RECT 107.900 39.600 109.700 39.900 ;
        RECT 107.900 39.500 108.200 39.600 ;
        RECT 105.400 36.600 105.700 36.900 ;
        RECT 103.900 36.300 105.700 36.600 ;
        RECT 106.300 36.700 106.600 36.900 ;
        RECT 107.800 36.700 108.200 39.500 ;
        RECT 109.400 39.500 109.700 39.600 ;
        RECT 106.300 36.500 108.200 36.700 ;
        RECT 108.600 36.500 109.000 39.300 ;
        RECT 109.400 36.500 109.800 39.500 ;
        RECT 106.300 36.400 108.100 36.500 ;
        RECT 108.600 36.200 108.900 36.500 ;
        RECT 110.500 36.300 110.900 39.900 ;
        RECT 108.600 36.100 109.000 36.200 ;
        RECT 101.300 35.500 102.500 35.800 ;
        RECT 107.300 35.800 109.000 36.100 ;
        RECT 110.500 35.900 111.400 36.300 ;
        RECT 100.600 34.800 101.000 35.200 ;
        RECT 100.600 33.100 100.900 34.800 ;
        RECT 101.300 33.800 101.600 35.500 ;
        RECT 102.200 34.800 102.600 35.200 ;
        RECT 106.200 34.800 107.000 35.200 ;
        RECT 102.200 34.400 102.500 34.800 ;
        RECT 102.000 34.000 102.600 34.400 ;
        RECT 103.000 33.800 103.400 34.600 ;
        RECT 104.600 34.100 105.000 34.200 ;
        RECT 105.400 34.100 106.200 34.200 ;
        RECT 104.600 33.800 106.200 34.100 ;
        RECT 101.200 33.700 101.600 33.800 ;
        RECT 101.200 33.500 102.700 33.700 ;
        RECT 101.200 33.400 103.300 33.500 ;
        RECT 102.400 33.200 103.300 33.400 ;
        RECT 103.000 33.100 103.300 33.200 ;
        RECT 100.600 32.600 101.300 33.100 ;
        RECT 100.900 31.100 101.300 32.600 ;
        RECT 103.000 31.100 103.400 33.100 ;
        RECT 104.600 32.800 105.500 33.200 ;
        RECT 107.300 32.500 107.600 35.800 ;
        RECT 110.200 34.800 110.600 35.600 ;
        RECT 111.000 34.200 111.300 35.900 ;
        RECT 112.600 35.600 113.000 39.900 ;
        RECT 114.700 37.900 115.300 39.900 ;
        RECT 117.000 37.900 117.400 39.900 ;
        RECT 119.200 38.200 119.600 39.900 ;
        RECT 119.200 37.900 120.200 38.200 ;
        RECT 115.000 37.500 115.400 37.900 ;
        RECT 117.100 37.600 117.400 37.900 ;
        RECT 116.700 37.300 118.500 37.600 ;
        RECT 119.800 37.500 120.200 37.900 ;
        RECT 116.700 37.200 117.100 37.300 ;
        RECT 118.100 37.200 118.500 37.300 ;
        RECT 114.600 36.600 115.300 37.000 ;
        RECT 114.200 35.600 114.600 36.200 ;
        RECT 115.000 36.100 115.300 36.600 ;
        RECT 116.100 36.500 117.200 36.800 ;
        RECT 116.100 36.400 116.500 36.500 ;
        RECT 115.000 35.800 116.200 36.100 ;
        RECT 112.600 35.300 114.700 35.600 ;
        RECT 111.000 33.800 111.400 34.200 ;
        RECT 110.200 33.100 110.600 33.200 ;
        RECT 111.000 33.100 111.300 33.800 ;
        RECT 112.600 33.600 113.000 35.300 ;
        RECT 114.300 35.200 114.700 35.300 ;
        RECT 113.500 34.900 113.900 35.000 ;
        RECT 113.500 34.600 115.400 34.900 ;
        RECT 115.000 34.500 115.400 34.600 ;
        RECT 115.900 34.200 116.200 35.800 ;
        RECT 116.900 35.900 117.200 36.500 ;
        RECT 117.500 36.500 117.900 36.600 ;
        RECT 119.800 36.500 120.200 36.600 ;
        RECT 117.500 36.200 120.200 36.500 ;
        RECT 116.900 35.700 119.300 35.900 ;
        RECT 121.400 35.700 121.800 39.900 ;
        RECT 123.500 36.300 123.900 39.900 ;
        RECT 123.000 35.900 123.900 36.300 ;
        RECT 116.900 35.600 121.800 35.700 ;
        RECT 118.900 35.500 121.800 35.600 ;
        RECT 119.000 35.400 121.800 35.500 ;
        RECT 118.200 35.100 118.600 35.200 ;
        RECT 118.200 34.800 120.700 35.100 ;
        RECT 119.000 34.700 119.400 34.800 ;
        RECT 120.300 34.700 120.700 34.800 ;
        RECT 119.500 34.200 119.900 34.300 ;
        RECT 123.100 34.200 123.400 35.900 ;
        RECT 124.600 35.600 125.000 39.900 ;
        RECT 126.700 37.900 127.300 39.900 ;
        RECT 129.000 37.900 129.400 39.900 ;
        RECT 131.200 38.200 131.600 39.900 ;
        RECT 131.200 37.900 132.200 38.200 ;
        RECT 127.000 37.500 127.400 37.900 ;
        RECT 129.100 37.600 129.400 37.900 ;
        RECT 128.700 37.300 130.500 37.600 ;
        RECT 131.800 37.500 132.200 37.900 ;
        RECT 128.700 37.200 129.100 37.300 ;
        RECT 130.100 37.200 130.500 37.300 ;
        RECT 126.600 36.600 127.300 37.000 ;
        RECT 127.000 36.100 127.300 36.600 ;
        RECT 128.100 36.500 129.200 36.800 ;
        RECT 128.100 36.400 128.500 36.500 ;
        RECT 127.000 35.800 128.200 36.100 ;
        RECT 123.800 34.800 124.200 35.600 ;
        RECT 124.600 35.300 126.700 35.600 ;
        RECT 115.900 33.900 121.400 34.200 ;
        RECT 116.100 33.800 116.500 33.900 ;
        RECT 112.600 33.300 114.500 33.600 ;
        RECT 110.200 32.800 111.300 33.100 ;
        RECT 105.600 32.200 107.600 32.500 ;
        RECT 105.400 31.800 105.900 32.200 ;
        RECT 107.000 32.100 107.600 32.200 ;
        RECT 111.000 32.100 111.300 32.800 ;
        RECT 111.800 32.400 112.200 33.200 ;
        RECT 105.400 31.100 105.800 31.800 ;
        RECT 107.000 31.100 107.400 32.100 ;
        RECT 111.000 31.100 111.400 32.100 ;
        RECT 112.600 31.100 113.000 33.300 ;
        RECT 114.100 33.200 114.500 33.300 ;
        RECT 119.000 32.800 119.300 33.900 ;
        RECT 120.600 33.800 121.400 33.900 ;
        RECT 123.000 33.800 123.400 34.200 ;
        RECT 118.100 32.700 118.500 32.800 ;
        RECT 115.000 32.100 115.400 32.500 ;
        RECT 117.100 32.400 118.500 32.700 ;
        RECT 119.000 32.400 119.400 32.800 ;
        RECT 117.100 32.100 117.400 32.400 ;
        RECT 119.800 32.100 120.200 32.500 ;
        RECT 114.700 31.800 115.400 32.100 ;
        RECT 114.700 31.100 115.300 31.800 ;
        RECT 117.000 31.100 117.400 32.100 ;
        RECT 119.200 31.800 120.200 32.100 ;
        RECT 119.200 31.100 119.600 31.800 ;
        RECT 121.400 31.100 121.800 33.500 ;
        RECT 122.200 32.400 122.600 33.200 ;
        RECT 123.100 32.100 123.400 33.800 ;
        RECT 123.000 31.100 123.400 32.100 ;
        RECT 124.600 33.600 125.000 35.300 ;
        RECT 126.300 35.200 126.700 35.300 ;
        RECT 125.500 34.900 125.900 35.000 ;
        RECT 125.500 34.600 127.400 34.900 ;
        RECT 127.000 34.500 127.400 34.600 ;
        RECT 127.900 34.200 128.200 35.800 ;
        RECT 128.900 35.900 129.200 36.500 ;
        RECT 129.500 36.500 129.900 36.600 ;
        RECT 131.800 36.500 132.200 36.600 ;
        RECT 129.500 36.200 132.200 36.500 ;
        RECT 128.900 35.700 131.300 35.900 ;
        RECT 133.400 35.700 133.800 39.900 ;
        RECT 128.900 35.600 133.800 35.700 ;
        RECT 130.900 35.500 133.800 35.600 ;
        RECT 131.000 35.400 133.800 35.500 ;
        RECT 134.200 35.900 134.600 39.900 ;
        RECT 135.800 36.200 136.200 39.900 ;
        RECT 135.100 35.900 136.200 36.200 ;
        RECT 136.600 36.200 137.000 39.900 ;
        RECT 136.600 35.900 137.700 36.200 ;
        RECT 138.200 35.900 138.600 39.900 ;
        RECT 130.200 35.100 130.600 35.200 ;
        RECT 130.200 34.800 132.700 35.100 ;
        RECT 132.300 34.700 132.700 34.800 ;
        RECT 134.200 34.800 134.500 35.900 ;
        RECT 135.100 35.600 135.400 35.900 ;
        RECT 134.800 35.200 135.400 35.600 ;
        RECT 131.500 34.200 131.900 34.300 ;
        RECT 127.900 33.900 133.400 34.200 ;
        RECT 128.100 33.800 128.500 33.900 ;
        RECT 129.400 33.800 129.800 33.900 ;
        RECT 124.600 33.300 126.500 33.600 ;
        RECT 124.600 31.100 125.000 33.300 ;
        RECT 126.100 33.200 126.500 33.300 ;
        RECT 131.000 32.800 131.300 33.900 ;
        RECT 132.600 33.800 133.400 33.900 ;
        RECT 130.100 32.700 130.500 32.800 ;
        RECT 127.000 32.100 127.400 32.500 ;
        RECT 129.100 32.400 130.500 32.700 ;
        RECT 131.000 32.400 131.400 32.800 ;
        RECT 129.100 32.100 129.400 32.400 ;
        RECT 131.800 32.100 132.200 32.500 ;
        RECT 126.700 31.800 127.400 32.100 ;
        RECT 126.700 31.100 127.300 31.800 ;
        RECT 129.000 31.100 129.400 32.100 ;
        RECT 131.200 31.800 132.200 32.100 ;
        RECT 131.200 31.100 131.600 31.800 ;
        RECT 133.400 31.100 133.800 33.500 ;
        RECT 134.200 31.100 134.600 34.800 ;
        RECT 135.100 33.700 135.400 35.200 ;
        RECT 137.400 35.600 137.700 35.900 ;
        RECT 137.400 35.200 138.000 35.600 ;
        RECT 137.400 33.700 137.700 35.200 ;
        RECT 138.300 34.800 138.600 35.900 ;
        RECT 139.800 35.600 140.200 39.900 ;
        RECT 141.400 35.600 141.800 39.900 ;
        RECT 143.000 35.600 143.400 39.900 ;
        RECT 144.600 35.600 145.000 39.900 ;
        RECT 147.800 35.700 148.200 39.900 ;
        RECT 150.000 38.200 150.400 39.900 ;
        RECT 149.400 37.900 150.400 38.200 ;
        RECT 152.200 37.900 152.600 39.900 ;
        RECT 154.300 37.900 154.900 39.900 ;
        RECT 149.400 37.500 149.800 37.900 ;
        RECT 152.200 37.600 152.500 37.900 ;
        RECT 151.100 37.300 152.900 37.600 ;
        RECT 154.200 37.500 154.600 37.900 ;
        RECT 151.100 37.200 151.500 37.300 ;
        RECT 152.500 37.200 152.900 37.300 ;
        RECT 149.400 36.500 149.800 36.600 ;
        RECT 151.700 36.500 152.100 36.600 ;
        RECT 149.400 36.200 152.100 36.500 ;
        RECT 152.400 36.500 153.500 36.800 ;
        RECT 152.400 35.900 152.700 36.500 ;
        RECT 153.100 36.400 153.500 36.500 ;
        RECT 154.300 36.600 155.000 37.000 ;
        RECT 154.300 36.100 154.600 36.600 ;
        RECT 150.300 35.700 152.700 35.900 ;
        RECT 147.800 35.600 152.700 35.700 ;
        RECT 153.400 35.800 154.600 36.100 ;
        RECT 139.800 35.200 140.700 35.600 ;
        RECT 141.400 35.200 142.500 35.600 ;
        RECT 143.000 35.200 144.100 35.600 ;
        RECT 144.600 35.200 145.800 35.600 ;
        RECT 147.800 35.500 150.700 35.600 ;
        RECT 147.800 35.400 150.600 35.500 ;
        RECT 135.100 33.400 136.200 33.700 ;
        RECT 135.800 31.100 136.200 33.400 ;
        RECT 136.600 33.400 137.700 33.700 ;
        RECT 136.600 31.100 137.000 33.400 ;
        RECT 138.200 31.100 138.600 34.800 ;
        RECT 140.300 34.500 140.700 35.200 ;
        RECT 142.100 34.500 142.500 35.200 ;
        RECT 143.700 34.500 144.100 35.200 ;
        RECT 140.300 34.100 141.600 34.500 ;
        RECT 142.100 34.100 143.300 34.500 ;
        RECT 143.700 34.100 145.000 34.500 ;
        RECT 140.300 33.800 140.700 34.100 ;
        RECT 142.100 33.800 142.500 34.100 ;
        RECT 143.700 33.800 144.100 34.100 ;
        RECT 145.400 33.800 145.800 35.200 ;
        RECT 151.000 35.100 151.400 35.200 ;
        RECT 148.900 34.800 151.400 35.100 ;
        RECT 148.900 34.700 149.300 34.800 ;
        RECT 149.700 34.200 150.100 34.300 ;
        RECT 153.400 34.200 153.700 35.800 ;
        RECT 156.600 35.600 157.000 39.900 ;
        RECT 154.900 35.300 157.000 35.600 ;
        RECT 157.400 35.700 157.800 39.900 ;
        RECT 159.600 38.200 160.000 39.900 ;
        RECT 159.000 37.900 160.000 38.200 ;
        RECT 161.800 37.900 162.200 39.900 ;
        RECT 163.900 37.900 164.500 39.900 ;
        RECT 159.000 37.500 159.400 37.900 ;
        RECT 161.800 37.600 162.100 37.900 ;
        RECT 160.700 37.300 162.500 37.600 ;
        RECT 163.800 37.500 164.200 37.900 ;
        RECT 160.700 37.200 161.100 37.300 ;
        RECT 162.100 37.200 162.500 37.300 ;
        RECT 159.000 36.500 159.400 36.600 ;
        RECT 161.300 36.500 161.700 36.600 ;
        RECT 159.000 36.200 161.700 36.500 ;
        RECT 162.000 36.500 163.100 36.800 ;
        RECT 162.000 35.900 162.300 36.500 ;
        RECT 162.700 36.400 163.100 36.500 ;
        RECT 163.900 36.600 164.600 37.000 ;
        RECT 163.900 36.100 164.200 36.600 ;
        RECT 159.900 35.700 162.300 35.900 ;
        RECT 157.400 35.600 162.300 35.700 ;
        RECT 163.000 35.800 164.200 36.100 ;
        RECT 157.400 35.500 160.300 35.600 ;
        RECT 157.400 35.400 160.200 35.500 ;
        RECT 154.900 35.200 155.300 35.300 ;
        RECT 155.700 34.900 156.100 35.000 ;
        RECT 154.200 34.600 156.100 34.900 ;
        RECT 154.200 34.500 154.600 34.600 ;
        RECT 148.200 33.900 153.700 34.200 ;
        RECT 148.200 33.800 149.000 33.900 ;
        RECT 139.800 33.400 140.700 33.800 ;
        RECT 141.400 33.400 142.500 33.800 ;
        RECT 143.000 33.400 144.100 33.800 ;
        RECT 144.600 33.400 145.800 33.800 ;
        RECT 139.800 31.100 140.200 33.400 ;
        RECT 141.400 31.100 141.800 33.400 ;
        RECT 143.000 31.100 143.400 33.400 ;
        RECT 144.600 31.100 145.000 33.400 ;
        RECT 147.800 31.100 148.200 33.500 ;
        RECT 150.300 33.200 150.600 33.900 ;
        RECT 153.100 33.800 153.500 33.900 ;
        RECT 156.600 33.600 157.000 35.300 ;
        RECT 160.600 35.100 161.000 35.200 ;
        RECT 162.200 35.100 162.600 35.200 ;
        RECT 158.500 34.800 162.600 35.100 ;
        RECT 158.500 34.700 158.900 34.800 ;
        RECT 159.300 34.200 159.700 34.300 ;
        RECT 163.000 34.200 163.300 35.800 ;
        RECT 166.200 35.600 166.600 39.900 ;
        RECT 167.000 35.900 167.400 39.900 ;
        RECT 167.800 36.200 168.200 39.900 ;
        RECT 169.400 36.200 169.800 39.900 ;
        RECT 167.800 35.900 169.800 36.200 ;
        RECT 164.500 35.300 166.600 35.600 ;
        RECT 164.500 35.200 164.900 35.300 ;
        RECT 165.300 34.900 165.700 35.000 ;
        RECT 163.800 34.600 165.700 34.900 ;
        RECT 163.800 34.500 164.200 34.600 ;
        RECT 157.800 33.900 163.300 34.200 ;
        RECT 157.800 33.800 158.600 33.900 ;
        RECT 155.100 33.300 157.000 33.600 ;
        RECT 155.100 33.200 155.500 33.300 ;
        RECT 149.400 32.100 149.800 32.500 ;
        RECT 150.200 32.400 150.600 33.200 ;
        RECT 151.100 32.700 151.500 32.800 ;
        RECT 151.100 32.400 152.500 32.700 ;
        RECT 152.200 32.100 152.500 32.400 ;
        RECT 154.200 32.100 154.600 32.500 ;
        RECT 149.400 31.800 150.400 32.100 ;
        RECT 150.000 31.100 150.400 31.800 ;
        RECT 152.200 31.100 152.600 32.100 ;
        RECT 154.200 31.800 154.900 32.100 ;
        RECT 154.300 31.100 154.900 31.800 ;
        RECT 156.600 31.100 157.000 33.300 ;
        RECT 157.400 31.100 157.800 33.500 ;
        RECT 159.900 32.800 160.200 33.900 ;
        RECT 162.700 33.800 163.100 33.900 ;
        RECT 166.200 33.600 166.600 35.300 ;
        RECT 167.100 35.200 167.400 35.900 ;
        RECT 170.200 35.600 170.600 39.900 ;
        RECT 172.300 37.900 172.900 39.900 ;
        RECT 174.600 37.900 175.000 39.900 ;
        RECT 176.800 38.200 177.200 39.900 ;
        RECT 176.800 37.900 177.800 38.200 ;
        RECT 172.600 37.500 173.000 37.900 ;
        RECT 174.700 37.600 175.000 37.900 ;
        RECT 174.300 37.300 176.100 37.600 ;
        RECT 177.400 37.500 177.800 37.900 ;
        RECT 174.300 37.200 174.700 37.300 ;
        RECT 175.700 37.200 176.100 37.300 ;
        RECT 172.200 36.600 172.900 37.000 ;
        RECT 172.600 36.100 172.900 36.600 ;
        RECT 173.700 36.500 174.800 36.800 ;
        RECT 173.700 36.400 174.100 36.500 ;
        RECT 172.600 35.800 173.800 36.100 ;
        RECT 169.000 35.200 169.400 35.400 ;
        RECT 170.200 35.300 172.300 35.600 ;
        RECT 167.000 34.900 168.200 35.200 ;
        RECT 169.000 35.100 169.800 35.200 ;
        RECT 170.200 35.100 170.600 35.300 ;
        RECT 171.900 35.200 172.300 35.300 ;
        RECT 173.500 35.200 173.800 35.800 ;
        RECT 174.500 35.900 174.800 36.500 ;
        RECT 175.100 36.500 175.500 36.600 ;
        RECT 177.400 36.500 177.800 36.600 ;
        RECT 175.100 36.200 177.800 36.500 ;
        RECT 174.500 35.700 176.900 35.900 ;
        RECT 179.000 35.700 179.400 39.900 ;
        RECT 174.500 35.600 179.400 35.700 ;
        RECT 176.500 35.500 179.400 35.600 ;
        RECT 176.600 35.400 179.400 35.500 ;
        RECT 179.800 35.700 180.200 39.900 ;
        RECT 182.000 38.200 182.400 39.900 ;
        RECT 181.400 37.900 182.400 38.200 ;
        RECT 184.200 37.900 184.600 39.900 ;
        RECT 186.300 37.900 186.900 39.900 ;
        RECT 181.400 37.500 181.800 37.900 ;
        RECT 184.200 37.600 184.500 37.900 ;
        RECT 183.100 37.300 184.900 37.600 ;
        RECT 186.200 37.500 186.600 37.900 ;
        RECT 183.100 37.200 183.500 37.300 ;
        RECT 184.500 37.200 184.900 37.300 ;
        RECT 186.700 37.000 187.400 37.200 ;
        RECT 186.300 36.800 187.400 37.000 ;
        RECT 181.400 36.500 181.800 36.600 ;
        RECT 183.700 36.500 184.100 36.600 ;
        RECT 181.400 36.200 184.100 36.500 ;
        RECT 184.400 36.500 185.500 36.800 ;
        RECT 184.400 35.900 184.700 36.500 ;
        RECT 185.100 36.400 185.500 36.500 ;
        RECT 186.300 36.600 187.000 36.800 ;
        RECT 186.300 36.100 186.600 36.600 ;
        RECT 182.300 35.700 184.700 35.900 ;
        RECT 179.800 35.600 184.700 35.700 ;
        RECT 185.400 35.800 186.600 36.100 ;
        RECT 179.800 35.500 182.700 35.600 ;
        RECT 179.800 35.400 182.600 35.500 ;
        RECT 169.000 34.900 170.600 35.100 ;
        RECT 167.000 34.800 167.400 34.900 ;
        RECT 167.800 34.800 168.200 34.900 ;
        RECT 169.400 34.800 170.600 34.900 ;
        RECT 164.700 33.300 166.600 33.600 ;
        RECT 164.700 33.200 165.100 33.300 ;
        RECT 159.000 32.100 159.400 32.500 ;
        RECT 159.800 32.400 160.200 32.800 ;
        RECT 160.700 32.700 161.100 32.800 ;
        RECT 160.700 32.400 162.100 32.700 ;
        RECT 161.800 32.100 162.100 32.400 ;
        RECT 163.800 32.100 164.200 32.500 ;
        RECT 159.000 31.800 160.000 32.100 ;
        RECT 159.600 31.100 160.000 31.800 ;
        RECT 161.800 31.100 162.200 32.100 ;
        RECT 163.800 31.800 164.500 32.100 ;
        RECT 163.900 31.100 164.500 31.800 ;
        RECT 166.200 31.100 166.600 33.300 ;
        RECT 167.000 32.800 167.400 33.200 ;
        RECT 167.900 33.100 168.200 34.800 ;
        RECT 168.600 33.800 169.000 34.600 ;
        RECT 167.100 32.400 167.500 32.800 ;
        RECT 167.800 31.100 168.200 33.100 ;
        RECT 170.200 33.600 170.600 34.800 ;
        RECT 171.100 34.900 171.500 35.000 ;
        RECT 171.100 34.600 173.000 34.900 ;
        RECT 173.400 34.800 173.800 35.200 ;
        RECT 175.800 35.100 176.200 35.200 ;
        RECT 183.000 35.100 183.400 35.200 ;
        RECT 175.800 34.800 178.300 35.100 ;
        RECT 172.600 34.500 173.000 34.600 ;
        RECT 173.500 34.200 173.800 34.800 ;
        RECT 177.900 34.700 178.300 34.800 ;
        RECT 180.900 34.800 183.400 35.100 ;
        RECT 180.900 34.700 181.300 34.800 ;
        RECT 182.200 34.700 182.600 34.800 ;
        RECT 177.100 34.200 177.500 34.300 ;
        RECT 181.700 34.200 182.100 34.300 ;
        RECT 185.400 34.200 185.700 35.800 ;
        RECT 188.600 35.600 189.000 39.900 ;
        RECT 189.400 36.200 189.800 39.900 ;
        RECT 189.400 35.900 190.500 36.200 ;
        RECT 191.000 35.900 191.400 39.900 ;
        RECT 191.800 36.200 192.200 39.900 ;
        RECT 191.800 35.900 192.900 36.200 ;
        RECT 193.400 35.900 193.800 39.900 ;
        RECT 186.900 35.300 189.000 35.600 ;
        RECT 186.900 35.200 187.300 35.300 ;
        RECT 187.700 34.900 188.100 35.000 ;
        RECT 186.200 34.600 188.100 34.900 ;
        RECT 186.200 34.500 186.600 34.600 ;
        RECT 173.500 34.100 179.000 34.200 ;
        RECT 180.200 34.100 185.700 34.200 ;
        RECT 173.500 33.900 185.700 34.100 ;
        RECT 173.700 33.800 174.100 33.900 ;
        RECT 170.200 33.300 172.100 33.600 ;
        RECT 170.200 31.100 170.600 33.300 ;
        RECT 171.700 33.200 172.100 33.300 ;
        RECT 176.600 32.800 176.900 33.900 ;
        RECT 178.200 33.800 181.000 33.900 ;
        RECT 175.700 32.700 176.100 32.800 ;
        RECT 172.600 32.100 173.000 32.500 ;
        RECT 174.700 32.400 176.100 32.700 ;
        RECT 176.600 32.400 177.000 32.800 ;
        RECT 174.700 32.100 175.000 32.400 ;
        RECT 177.400 32.100 177.800 32.500 ;
        RECT 172.300 31.800 173.000 32.100 ;
        RECT 172.300 31.100 172.900 31.800 ;
        RECT 174.600 31.100 175.000 32.100 ;
        RECT 176.800 31.800 177.800 32.100 ;
        RECT 176.800 31.100 177.200 31.800 ;
        RECT 179.000 31.100 179.400 33.500 ;
        RECT 179.800 31.100 180.200 33.500 ;
        RECT 182.300 32.800 182.600 33.900 ;
        RECT 185.100 33.800 185.500 33.900 ;
        RECT 188.600 33.600 189.000 35.300 ;
        RECT 190.200 35.600 190.500 35.900 ;
        RECT 190.200 35.200 190.800 35.600 ;
        RECT 190.200 33.700 190.500 35.200 ;
        RECT 191.100 34.800 191.400 35.900 ;
        RECT 187.100 33.300 189.000 33.600 ;
        RECT 187.100 33.200 187.500 33.300 ;
        RECT 181.400 32.100 181.800 32.500 ;
        RECT 182.200 32.400 182.600 32.800 ;
        RECT 183.100 32.700 183.500 32.800 ;
        RECT 183.100 32.400 184.500 32.700 ;
        RECT 184.200 32.100 184.500 32.400 ;
        RECT 186.200 32.100 186.600 32.500 ;
        RECT 181.400 31.800 182.400 32.100 ;
        RECT 182.000 31.100 182.400 31.800 ;
        RECT 184.200 31.100 184.600 32.100 ;
        RECT 186.200 31.800 186.900 32.100 ;
        RECT 186.300 31.100 186.900 31.800 ;
        RECT 188.600 31.100 189.000 33.300 ;
        RECT 189.400 33.400 190.500 33.700 ;
        RECT 189.400 31.100 189.800 33.400 ;
        RECT 191.000 31.100 191.400 34.800 ;
        RECT 192.600 35.600 192.900 35.900 ;
        RECT 192.600 35.200 193.200 35.600 ;
        RECT 192.600 33.700 192.900 35.200 ;
        RECT 193.500 34.800 193.800 35.900 ;
        RECT 191.800 33.400 192.900 33.700 ;
        RECT 191.800 31.100 192.200 33.400 ;
        RECT 193.400 31.100 193.800 34.800 ;
        RECT 1.400 28.900 1.800 29.900 ;
        RECT 1.500 27.800 1.800 28.900 ;
        RECT 3.000 27.900 3.400 29.900 ;
        RECT 4.600 28.900 5.000 29.900 ;
        RECT 1.500 27.500 2.700 27.800 ;
        RECT 1.400 26.800 1.900 27.200 ;
        RECT 1.600 26.400 2.000 26.800 ;
        RECT 2.400 26.000 2.700 27.500 ;
        RECT 3.100 26.200 3.400 27.900 ;
        RECT 3.800 27.800 4.200 28.600 ;
        RECT 4.700 27.800 5.000 28.900 ;
        RECT 6.200 27.900 6.600 29.900 ;
        RECT 4.700 27.500 5.900 27.800 ;
        RECT 2.300 25.700 2.700 26.000 ;
        RECT 3.000 25.800 3.400 26.200 ;
        RECT 5.600 26.000 5.900 27.500 ;
        RECT 6.300 26.200 6.600 27.900 ;
        RECT 0.600 25.600 2.700 25.700 ;
        RECT 0.600 25.400 2.600 25.600 ;
        RECT 0.600 21.100 1.000 25.400 ;
        RECT 3.100 25.100 3.400 25.800 ;
        RECT 5.500 25.700 5.900 26.000 ;
        RECT 6.200 25.800 6.600 26.200 ;
        RECT 2.700 24.800 3.400 25.100 ;
        RECT 3.800 25.600 5.900 25.700 ;
        RECT 3.800 25.400 5.800 25.600 ;
        RECT 2.700 21.100 3.100 24.800 ;
        RECT 3.800 21.100 4.200 25.400 ;
        RECT 6.300 25.100 6.600 25.800 ;
        RECT 5.900 24.800 6.600 25.100 ;
        RECT 5.900 21.100 6.300 24.800 ;
        RECT 7.000 24.100 7.400 24.200 ;
        RECT 7.800 24.100 8.200 29.900 ;
        RECT 8.600 27.500 9.000 29.900 ;
        RECT 10.800 29.200 11.200 29.900 ;
        RECT 10.200 28.900 11.200 29.200 ;
        RECT 13.000 28.900 13.400 29.900 ;
        RECT 15.100 29.200 15.700 29.900 ;
        RECT 15.000 28.900 15.700 29.200 ;
        RECT 10.200 28.500 10.600 28.900 ;
        RECT 13.000 28.600 13.300 28.900 ;
        RECT 11.000 28.200 11.400 28.600 ;
        RECT 11.900 28.300 13.300 28.600 ;
        RECT 15.000 28.500 15.400 28.900 ;
        RECT 11.900 28.200 12.300 28.300 ;
        RECT 9.000 27.100 9.800 27.200 ;
        RECT 11.100 27.100 11.400 28.200 ;
        RECT 14.200 27.800 14.600 28.200 ;
        RECT 14.200 27.200 14.500 27.800 ;
        RECT 15.900 27.700 16.300 27.800 ;
        RECT 17.400 27.700 17.800 29.900 ;
        RECT 15.900 27.400 17.800 27.700 ;
        RECT 18.200 27.500 18.600 29.900 ;
        RECT 20.400 29.200 20.800 29.900 ;
        RECT 19.800 28.900 20.800 29.200 ;
        RECT 22.600 28.900 23.000 29.900 ;
        RECT 24.700 29.200 25.300 29.900 ;
        RECT 24.600 28.900 25.300 29.200 ;
        RECT 19.800 28.500 20.200 28.900 ;
        RECT 22.600 28.600 22.900 28.900 ;
        RECT 20.600 28.200 21.000 28.600 ;
        RECT 21.500 28.300 22.900 28.600 ;
        RECT 24.600 28.500 25.000 28.900 ;
        RECT 21.500 28.200 21.900 28.300 ;
        RECT 13.900 27.100 14.500 27.200 ;
        RECT 9.000 26.800 14.500 27.100 ;
        RECT 10.500 26.700 10.900 26.800 ;
        RECT 9.700 26.200 10.100 26.300 ;
        RECT 9.700 25.900 12.200 26.200 ;
        RECT 11.800 25.800 12.200 25.900 ;
        RECT 7.000 23.800 8.200 24.100 ;
        RECT 7.800 21.100 8.200 23.800 ;
        RECT 8.600 25.500 11.400 25.600 ;
        RECT 8.600 25.400 11.500 25.500 ;
        RECT 8.600 25.300 13.500 25.400 ;
        RECT 8.600 21.100 9.000 25.300 ;
        RECT 11.100 25.100 13.500 25.300 ;
        RECT 10.200 24.500 12.900 24.800 ;
        RECT 10.200 24.400 10.600 24.500 ;
        RECT 12.500 24.400 12.900 24.500 ;
        RECT 13.200 24.500 13.500 25.100 ;
        RECT 14.200 25.200 14.500 26.800 ;
        RECT 15.000 26.400 15.400 26.500 ;
        RECT 15.000 26.100 16.900 26.400 ;
        RECT 16.500 26.000 16.900 26.100 ;
        RECT 15.700 25.700 16.100 25.800 ;
        RECT 17.400 25.700 17.800 27.400 ;
        RECT 18.600 27.100 19.400 27.200 ;
        RECT 20.700 27.100 21.000 28.200 ;
        RECT 25.500 27.700 25.900 27.800 ;
        RECT 27.000 27.700 27.400 29.900 ;
        RECT 25.500 27.400 27.400 27.700 ;
        RECT 27.800 27.500 28.200 29.900 ;
        RECT 30.000 29.200 30.400 29.900 ;
        RECT 29.400 28.900 30.400 29.200 ;
        RECT 32.200 28.900 32.600 29.900 ;
        RECT 34.300 29.200 34.900 29.900 ;
        RECT 34.200 28.900 34.900 29.200 ;
        RECT 29.400 28.500 29.800 28.900 ;
        RECT 32.200 28.600 32.500 28.900 ;
        RECT 30.200 28.200 30.600 28.600 ;
        RECT 31.100 28.300 32.500 28.600 ;
        RECT 34.200 28.500 34.600 28.900 ;
        RECT 31.100 28.200 31.500 28.300 ;
        RECT 23.500 27.100 23.900 27.200 ;
        RECT 18.600 26.800 24.100 27.100 ;
        RECT 20.100 26.700 20.500 26.800 ;
        RECT 19.300 26.200 19.700 26.300 ;
        RECT 20.600 26.200 21.000 26.300 ;
        RECT 23.800 26.200 24.100 26.800 ;
        RECT 24.600 26.400 25.000 26.500 ;
        RECT 19.300 25.900 21.800 26.200 ;
        RECT 21.400 25.800 21.800 25.900 ;
        RECT 23.800 25.800 24.200 26.200 ;
        RECT 24.600 26.100 26.500 26.400 ;
        RECT 26.100 26.000 26.500 26.100 ;
        RECT 15.700 25.400 17.800 25.700 ;
        RECT 14.200 24.900 15.400 25.200 ;
        RECT 13.900 24.500 14.300 24.600 ;
        RECT 13.200 24.200 14.300 24.500 ;
        RECT 15.100 24.400 15.400 24.900 ;
        RECT 15.100 24.000 15.800 24.400 ;
        RECT 11.900 23.700 12.300 23.800 ;
        RECT 13.300 23.700 13.700 23.800 ;
        RECT 10.200 23.100 10.600 23.500 ;
        RECT 11.900 23.400 13.700 23.700 ;
        RECT 13.000 23.100 13.300 23.400 ;
        RECT 15.000 23.100 15.400 23.500 ;
        RECT 10.200 22.800 11.200 23.100 ;
        RECT 10.800 21.100 11.200 22.800 ;
        RECT 13.000 21.100 13.400 23.100 ;
        RECT 15.100 21.100 15.700 23.100 ;
        RECT 17.400 21.100 17.800 25.400 ;
        RECT 18.200 25.500 21.000 25.600 ;
        RECT 18.200 25.400 21.100 25.500 ;
        RECT 18.200 25.300 23.100 25.400 ;
        RECT 18.200 21.100 18.600 25.300 ;
        RECT 20.700 25.100 23.100 25.300 ;
        RECT 19.800 24.500 22.500 24.800 ;
        RECT 19.800 24.400 20.200 24.500 ;
        RECT 22.100 24.400 22.500 24.500 ;
        RECT 22.800 24.500 23.100 25.100 ;
        RECT 23.800 25.200 24.100 25.800 ;
        RECT 25.300 25.700 25.700 25.800 ;
        RECT 27.000 25.700 27.400 27.400 ;
        RECT 28.200 27.100 29.000 27.200 ;
        RECT 30.300 27.100 30.600 28.200 ;
        RECT 35.100 27.700 35.500 27.800 ;
        RECT 36.600 27.700 37.000 29.900 ;
        RECT 35.100 27.400 37.000 27.700 ;
        RECT 33.100 27.100 33.500 27.200 ;
        RECT 28.200 26.800 33.700 27.100 ;
        RECT 29.700 26.700 30.100 26.800 ;
        RECT 28.900 26.200 29.300 26.300 ;
        RECT 30.200 26.200 30.600 26.300 ;
        RECT 28.900 25.900 31.400 26.200 ;
        RECT 31.000 25.800 31.400 25.900 ;
        RECT 25.300 25.400 27.400 25.700 ;
        RECT 23.800 24.900 25.000 25.200 ;
        RECT 23.500 24.500 23.900 24.600 ;
        RECT 22.800 24.200 23.900 24.500 ;
        RECT 24.700 24.400 25.000 24.900 ;
        RECT 24.700 24.000 25.400 24.400 ;
        RECT 21.500 23.700 21.900 23.800 ;
        RECT 22.900 23.700 23.300 23.800 ;
        RECT 19.800 23.100 20.200 23.500 ;
        RECT 21.500 23.400 23.300 23.700 ;
        RECT 22.600 23.100 22.900 23.400 ;
        RECT 24.600 23.100 25.000 23.500 ;
        RECT 19.800 22.800 20.800 23.100 ;
        RECT 20.400 21.100 20.800 22.800 ;
        RECT 22.600 21.100 23.000 23.100 ;
        RECT 24.700 21.100 25.300 23.100 ;
        RECT 27.000 21.100 27.400 25.400 ;
        RECT 27.800 25.500 30.600 25.600 ;
        RECT 27.800 25.400 30.700 25.500 ;
        RECT 27.800 25.300 32.700 25.400 ;
        RECT 27.800 21.100 28.200 25.300 ;
        RECT 30.300 25.100 32.700 25.300 ;
        RECT 29.400 24.500 32.100 24.800 ;
        RECT 29.400 24.400 29.800 24.500 ;
        RECT 31.700 24.400 32.100 24.500 ;
        RECT 32.400 24.500 32.700 25.100 ;
        RECT 33.400 25.200 33.700 26.800 ;
        RECT 34.200 26.400 34.600 26.500 ;
        RECT 34.200 26.100 36.100 26.400 ;
        RECT 35.700 26.000 36.100 26.100 ;
        RECT 34.900 25.700 35.300 25.800 ;
        RECT 36.600 25.700 37.000 27.400 ;
        RECT 38.200 28.800 38.600 29.900 ;
        RECT 38.200 27.200 38.500 28.800 ;
        RECT 39.000 27.800 39.400 28.600 ;
        RECT 39.800 27.500 40.200 29.900 ;
        RECT 42.000 29.200 42.400 29.900 ;
        RECT 41.400 28.900 42.400 29.200 ;
        RECT 44.200 28.900 44.600 29.900 ;
        RECT 46.300 29.200 46.900 29.900 ;
        RECT 46.200 28.900 46.900 29.200 ;
        RECT 41.400 28.500 41.800 28.900 ;
        RECT 44.200 28.600 44.500 28.900 ;
        RECT 42.200 28.200 42.600 28.600 ;
        RECT 43.100 28.300 44.500 28.600 ;
        RECT 46.200 28.500 46.600 28.900 ;
        RECT 43.100 28.200 43.500 28.300 ;
        RECT 38.200 26.800 38.600 27.200 ;
        RECT 40.200 27.100 41.000 27.200 ;
        RECT 42.300 27.100 42.600 28.200 ;
        RECT 47.100 27.700 47.500 27.800 ;
        RECT 48.600 27.700 49.000 29.900 ;
        RECT 51.000 27.900 51.400 29.900 ;
        RECT 53.100 28.400 53.500 29.900 ;
        RECT 53.100 27.900 53.800 28.400 ;
        RECT 47.100 27.400 49.000 27.700 ;
        RECT 51.100 27.800 51.400 27.900 ;
        RECT 51.100 27.600 52.000 27.800 ;
        RECT 51.100 27.500 53.200 27.600 ;
        RECT 45.100 27.100 45.500 27.200 ;
        RECT 40.200 26.800 45.700 27.100 ;
        RECT 34.900 25.400 37.000 25.700 ;
        RECT 37.400 25.400 37.800 26.200 ;
        RECT 33.400 24.900 34.600 25.200 ;
        RECT 33.100 24.500 33.500 24.600 ;
        RECT 32.400 24.200 33.500 24.500 ;
        RECT 34.300 24.400 34.600 24.900 ;
        RECT 34.300 24.000 35.000 24.400 ;
        RECT 31.100 23.700 31.500 23.800 ;
        RECT 32.500 23.700 32.900 23.800 ;
        RECT 29.400 23.100 29.800 23.500 ;
        RECT 31.100 23.400 32.900 23.700 ;
        RECT 32.200 23.100 32.500 23.400 ;
        RECT 34.200 23.100 34.600 23.500 ;
        RECT 29.400 22.800 30.400 23.100 ;
        RECT 30.000 21.100 30.400 22.800 ;
        RECT 32.200 21.100 32.600 23.100 ;
        RECT 34.300 21.100 34.900 23.100 ;
        RECT 36.600 21.100 37.000 25.400 ;
        RECT 38.200 25.100 38.500 26.800 ;
        RECT 41.700 26.700 42.100 26.800 ;
        RECT 40.900 26.200 41.300 26.300 ;
        RECT 42.200 26.200 42.600 26.300 ;
        RECT 40.900 25.900 43.400 26.200 ;
        RECT 43.000 25.800 43.400 25.900 ;
        RECT 39.800 25.500 42.600 25.600 ;
        RECT 39.800 25.400 42.700 25.500 ;
        RECT 39.800 25.300 44.700 25.400 ;
        RECT 37.700 24.700 38.600 25.100 ;
        RECT 37.700 21.100 38.100 24.700 ;
        RECT 39.800 21.100 40.200 25.300 ;
        RECT 42.300 25.100 44.700 25.300 ;
        RECT 41.400 24.500 44.100 24.800 ;
        RECT 41.400 24.400 41.800 24.500 ;
        RECT 43.700 24.400 44.100 24.500 ;
        RECT 44.400 24.500 44.700 25.100 ;
        RECT 45.400 25.200 45.700 26.800 ;
        RECT 46.200 26.400 46.600 26.500 ;
        RECT 46.200 26.100 48.100 26.400 ;
        RECT 47.700 26.000 48.100 26.100 ;
        RECT 46.900 25.700 47.300 25.800 ;
        RECT 48.600 25.700 49.000 27.400 ;
        RECT 51.700 27.300 53.200 27.500 ;
        RECT 52.800 27.200 53.200 27.300 ;
        RECT 51.000 26.400 51.400 27.200 ;
        RECT 52.000 26.900 52.400 27.000 ;
        RECT 51.900 26.600 52.400 26.900 ;
        RECT 51.900 26.200 52.200 26.600 ;
        RECT 51.800 25.800 52.200 26.200 ;
        RECT 46.900 25.400 49.000 25.700 ;
        RECT 52.800 25.500 53.100 27.200 ;
        RECT 53.500 26.200 53.800 27.900 ;
        RECT 53.400 25.800 53.800 26.200 ;
        RECT 45.400 24.900 46.600 25.200 ;
        RECT 45.100 24.500 45.500 24.600 ;
        RECT 44.400 24.200 45.500 24.500 ;
        RECT 46.300 24.400 46.600 24.900 ;
        RECT 46.300 24.000 47.000 24.400 ;
        RECT 43.100 23.700 43.500 23.800 ;
        RECT 44.500 23.700 44.900 23.800 ;
        RECT 41.400 23.100 41.800 23.500 ;
        RECT 43.100 23.400 44.900 23.700 ;
        RECT 44.200 23.100 44.500 23.400 ;
        RECT 46.200 23.100 46.600 23.500 ;
        RECT 41.400 22.800 42.400 23.100 ;
        RECT 42.000 21.100 42.400 22.800 ;
        RECT 44.200 21.100 44.600 23.100 ;
        RECT 46.300 21.100 46.900 23.100 ;
        RECT 48.600 21.100 49.000 25.400 ;
        RECT 51.900 25.200 53.100 25.500 ;
        RECT 51.900 23.100 52.200 25.200 ;
        RECT 53.500 25.100 53.800 25.800 ;
        RECT 51.800 21.100 52.200 23.100 ;
        RECT 53.400 21.100 53.800 25.100 ;
        RECT 54.200 27.700 54.600 29.900 ;
        RECT 56.300 29.200 56.900 29.900 ;
        RECT 56.300 28.900 57.000 29.200 ;
        RECT 58.600 28.900 59.000 29.900 ;
        RECT 60.800 29.200 61.200 29.900 ;
        RECT 60.800 28.900 61.800 29.200 ;
        RECT 56.600 28.500 57.000 28.900 ;
        RECT 58.700 28.600 59.000 28.900 ;
        RECT 58.700 28.300 60.100 28.600 ;
        RECT 59.700 28.200 60.100 28.300 ;
        RECT 60.600 28.200 61.000 28.600 ;
        RECT 61.400 28.500 61.800 28.900 ;
        RECT 55.700 27.700 56.100 27.800 ;
        RECT 54.200 27.400 56.100 27.700 ;
        RECT 54.200 25.700 54.600 27.400 ;
        RECT 57.700 27.100 58.100 27.200 ;
        RECT 59.800 27.100 60.200 27.200 ;
        RECT 60.600 27.100 60.900 28.200 ;
        RECT 63.000 27.500 63.400 29.900 ;
        RECT 62.200 27.100 63.000 27.200 ;
        RECT 57.500 26.800 63.000 27.100 ;
        RECT 56.600 26.400 57.000 26.500 ;
        RECT 55.100 26.100 57.000 26.400 ;
        RECT 55.100 26.000 55.500 26.100 ;
        RECT 55.900 25.700 56.300 25.800 ;
        RECT 54.200 25.400 56.300 25.700 ;
        RECT 54.200 21.100 54.600 25.400 ;
        RECT 57.500 25.200 57.800 26.800 ;
        RECT 61.100 26.700 61.500 26.800 ;
        RECT 60.600 26.200 61.000 26.300 ;
        RECT 61.900 26.200 62.300 26.300 ;
        RECT 59.800 25.900 62.300 26.200 ;
        RECT 63.800 26.200 64.200 29.900 ;
        RECT 65.400 27.600 65.800 29.900 ;
        RECT 64.700 27.300 65.800 27.600 ;
        RECT 66.200 27.900 66.600 29.900 ;
        RECT 67.800 28.900 68.200 29.900 ;
        RECT 70.200 28.900 70.600 29.900 ;
        RECT 59.800 25.800 60.200 25.900 ;
        RECT 60.600 25.500 63.400 25.600 ;
        RECT 60.500 25.400 63.400 25.500 ;
        RECT 56.600 24.900 57.800 25.200 ;
        RECT 58.500 25.300 63.400 25.400 ;
        RECT 58.500 25.100 60.900 25.300 ;
        RECT 56.600 24.400 56.900 24.900 ;
        RECT 56.200 24.000 56.900 24.400 ;
        RECT 57.700 24.500 58.100 24.600 ;
        RECT 58.500 24.500 58.800 25.100 ;
        RECT 57.700 24.200 58.800 24.500 ;
        RECT 59.100 24.500 61.800 24.800 ;
        RECT 59.100 24.400 59.500 24.500 ;
        RECT 61.400 24.400 61.800 24.500 ;
        RECT 58.300 23.700 58.700 23.800 ;
        RECT 59.700 23.700 60.100 23.800 ;
        RECT 56.600 23.100 57.000 23.500 ;
        RECT 58.300 23.400 60.100 23.700 ;
        RECT 58.700 23.100 59.000 23.400 ;
        RECT 61.400 23.100 61.800 23.500 ;
        RECT 56.300 21.100 56.900 23.100 ;
        RECT 58.600 21.100 59.000 23.100 ;
        RECT 60.800 22.800 61.800 23.100 ;
        RECT 60.800 21.100 61.200 22.800 ;
        RECT 63.000 21.100 63.400 25.300 ;
        RECT 63.800 25.100 64.100 26.200 ;
        RECT 64.700 25.800 65.000 27.300 ;
        RECT 65.400 25.800 65.800 26.600 ;
        RECT 66.200 26.200 66.500 27.900 ;
        RECT 67.800 27.800 68.100 28.900 ;
        RECT 69.400 27.800 69.800 28.600 ;
        RECT 66.900 27.500 68.100 27.800 ;
        RECT 66.200 25.800 66.600 26.200 ;
        RECT 66.900 26.000 67.200 27.500 ;
        RECT 70.300 27.200 70.600 28.900 ;
        RECT 71.800 27.800 72.200 28.600 ;
        RECT 67.700 26.800 68.200 27.200 ;
        RECT 70.200 26.800 70.600 27.200 ;
        RECT 67.600 26.400 68.000 26.800 ;
        RECT 64.400 25.400 65.000 25.800 ;
        RECT 64.700 25.100 65.000 25.400 ;
        RECT 66.200 25.100 66.500 25.800 ;
        RECT 66.900 25.700 67.300 26.000 ;
        RECT 66.900 25.600 69.000 25.700 ;
        RECT 67.000 25.400 69.000 25.600 ;
        RECT 63.800 21.100 64.200 25.100 ;
        RECT 64.700 24.800 65.800 25.100 ;
        RECT 66.200 24.800 66.900 25.100 ;
        RECT 65.400 21.100 65.800 24.800 ;
        RECT 66.500 21.100 66.900 24.800 ;
        RECT 68.600 21.100 69.000 25.400 ;
        RECT 70.300 25.100 70.600 26.800 ;
        RECT 71.000 26.100 71.400 26.200 ;
        RECT 71.800 26.100 72.200 26.200 ;
        RECT 71.000 25.800 72.200 26.100 ;
        RECT 71.000 25.400 71.400 25.800 ;
        RECT 70.200 24.700 71.100 25.100 ;
        RECT 70.700 21.100 71.100 24.700 ;
        RECT 72.600 21.100 73.000 29.900 ;
        RECT 75.200 27.100 75.600 29.900 ;
        RECT 75.200 26.900 76.100 27.100 ;
        RECT 75.300 26.800 76.100 26.900 ;
        RECT 74.200 25.800 75.000 26.200 ;
        RECT 73.400 24.800 73.800 25.600 ;
        RECT 75.800 25.200 76.100 26.800 ;
        RECT 76.600 26.100 77.000 26.200 ;
        RECT 77.400 26.100 77.800 29.900 ;
        RECT 76.600 25.800 77.800 26.100 ;
        RECT 75.800 24.800 76.200 25.200 ;
        RECT 74.200 23.800 74.600 24.200 ;
        RECT 75.000 23.800 75.400 24.600 ;
        RECT 74.200 23.500 74.500 23.800 ;
        RECT 75.800 23.500 76.100 24.800 ;
        RECT 74.200 23.200 76.100 23.500 ;
        RECT 74.200 21.100 74.600 23.200 ;
        RECT 75.800 23.100 76.100 23.200 ;
        RECT 75.800 21.100 76.200 23.100 ;
        RECT 77.400 21.100 77.800 25.800 ;
        RECT 78.200 27.700 78.600 29.900 ;
        RECT 80.300 29.200 80.900 29.900 ;
        RECT 80.300 28.900 81.000 29.200 ;
        RECT 82.600 28.900 83.000 29.900 ;
        RECT 84.800 29.200 85.200 29.900 ;
        RECT 84.800 28.900 85.800 29.200 ;
        RECT 80.600 28.500 81.000 28.900 ;
        RECT 82.700 28.600 83.000 28.900 ;
        RECT 82.700 28.300 84.100 28.600 ;
        RECT 83.700 28.200 84.100 28.300 ;
        RECT 84.600 28.200 85.000 28.600 ;
        RECT 85.400 28.500 85.800 28.900 ;
        RECT 79.700 27.700 80.100 27.800 ;
        RECT 78.200 27.400 80.100 27.700 ;
        RECT 78.200 25.700 78.600 27.400 ;
        RECT 81.700 27.100 82.100 27.200 ;
        RECT 83.800 27.100 84.200 27.200 ;
        RECT 84.600 27.100 84.900 28.200 ;
        RECT 87.000 27.500 87.400 29.900 ;
        RECT 87.800 27.700 88.200 29.900 ;
        RECT 89.900 29.200 90.500 29.900 ;
        RECT 89.900 28.900 90.600 29.200 ;
        RECT 92.200 28.900 92.600 29.900 ;
        RECT 94.400 29.200 94.800 29.900 ;
        RECT 94.400 28.900 95.400 29.200 ;
        RECT 90.200 28.500 90.600 28.900 ;
        RECT 92.300 28.600 92.600 28.900 ;
        RECT 92.300 28.300 93.700 28.600 ;
        RECT 93.300 28.200 93.700 28.300 ;
        RECT 94.200 28.200 94.600 28.600 ;
        RECT 95.000 28.500 95.400 28.900 ;
        RECT 89.300 27.700 89.700 27.800 ;
        RECT 87.800 27.400 89.700 27.700 ;
        RECT 86.200 27.100 87.000 27.200 ;
        RECT 81.500 26.800 87.000 27.100 ;
        RECT 80.600 26.400 81.000 26.500 ;
        RECT 79.100 26.100 81.000 26.400 ;
        RECT 79.100 26.000 79.500 26.100 ;
        RECT 79.900 25.700 80.300 25.800 ;
        RECT 78.200 25.400 80.300 25.700 ;
        RECT 78.200 21.100 78.600 25.400 ;
        RECT 81.500 25.200 81.800 26.800 ;
        RECT 85.100 26.700 85.500 26.800 ;
        RECT 84.600 26.200 85.000 26.300 ;
        RECT 85.900 26.200 86.300 26.300 ;
        RECT 83.800 25.900 86.300 26.200 ;
        RECT 83.800 25.800 84.200 25.900 ;
        RECT 87.800 25.700 88.200 27.400 ;
        RECT 91.300 27.100 92.200 27.200 ;
        RECT 94.200 27.100 94.500 28.200 ;
        RECT 96.600 27.500 97.000 29.900 ;
        RECT 99.000 27.900 99.400 29.900 ;
        RECT 101.100 28.400 101.500 29.900 ;
        RECT 101.100 27.900 101.800 28.400 ;
        RECT 99.100 27.800 99.400 27.900 ;
        RECT 99.100 27.600 100.000 27.800 ;
        RECT 99.100 27.500 101.200 27.600 ;
        RECT 99.700 27.300 101.200 27.500 ;
        RECT 100.800 27.200 101.200 27.300 ;
        RECT 95.800 27.100 96.600 27.200 ;
        RECT 91.100 26.800 96.600 27.100 ;
        RECT 90.200 26.400 90.600 26.500 ;
        RECT 88.700 26.100 90.600 26.400 ;
        RECT 88.700 26.000 89.100 26.100 ;
        RECT 89.500 25.700 89.900 25.800 ;
        RECT 84.600 25.500 87.400 25.600 ;
        RECT 84.500 25.400 87.400 25.500 ;
        RECT 80.600 24.900 81.800 25.200 ;
        RECT 82.500 25.300 87.400 25.400 ;
        RECT 82.500 25.100 84.900 25.300 ;
        RECT 80.600 24.400 80.900 24.900 ;
        RECT 80.200 24.000 80.900 24.400 ;
        RECT 81.700 24.500 82.100 24.600 ;
        RECT 82.500 24.500 82.800 25.100 ;
        RECT 81.700 24.200 82.800 24.500 ;
        RECT 83.100 24.500 85.800 24.800 ;
        RECT 83.100 24.400 83.500 24.500 ;
        RECT 85.400 24.400 85.800 24.500 ;
        RECT 82.300 23.700 82.700 23.800 ;
        RECT 83.700 23.700 84.100 23.800 ;
        RECT 80.600 23.100 81.000 23.500 ;
        RECT 82.300 23.400 84.100 23.700 ;
        RECT 82.700 23.100 83.000 23.400 ;
        RECT 85.400 23.100 85.800 23.500 ;
        RECT 80.300 21.100 80.900 23.100 ;
        RECT 82.600 21.100 83.000 23.100 ;
        RECT 84.800 22.800 85.800 23.100 ;
        RECT 84.800 21.100 85.200 22.800 ;
        RECT 87.000 21.100 87.400 25.300 ;
        RECT 87.800 25.400 89.900 25.700 ;
        RECT 87.800 21.100 88.200 25.400 ;
        RECT 91.100 25.200 91.400 26.800 ;
        RECT 94.700 26.700 95.100 26.800 ;
        RECT 99.000 26.400 99.400 27.200 ;
        RECT 100.000 26.900 100.400 27.000 ;
        RECT 99.900 26.600 100.400 26.900 ;
        RECT 95.500 26.200 95.900 26.300 ;
        RECT 99.900 26.200 100.200 26.600 ;
        RECT 93.400 25.900 95.900 26.200 ;
        RECT 93.400 25.800 93.800 25.900 ;
        RECT 99.800 25.800 100.200 26.200 ;
        RECT 94.200 25.500 97.000 25.600 ;
        RECT 100.800 25.500 101.100 27.200 ;
        RECT 101.500 26.200 101.800 27.900 ;
        RECT 101.400 25.800 101.800 26.200 ;
        RECT 94.100 25.400 97.000 25.500 ;
        RECT 90.200 24.900 91.400 25.200 ;
        RECT 92.100 25.300 97.000 25.400 ;
        RECT 92.100 25.100 94.500 25.300 ;
        RECT 90.200 24.400 90.500 24.900 ;
        RECT 89.800 24.000 90.500 24.400 ;
        RECT 91.300 24.500 91.700 24.600 ;
        RECT 92.100 24.500 92.400 25.100 ;
        RECT 91.300 24.200 92.400 24.500 ;
        RECT 92.700 24.500 95.400 24.800 ;
        RECT 92.700 24.400 93.100 24.500 ;
        RECT 95.000 24.400 95.400 24.500 ;
        RECT 91.900 23.700 92.300 23.800 ;
        RECT 93.300 23.700 93.700 23.800 ;
        RECT 90.200 23.100 90.600 23.500 ;
        RECT 91.900 23.400 93.700 23.700 ;
        RECT 92.300 23.100 92.600 23.400 ;
        RECT 95.000 23.100 95.400 23.500 ;
        RECT 89.900 21.100 90.500 23.100 ;
        RECT 92.200 21.100 92.600 23.100 ;
        RECT 94.400 22.800 95.400 23.100 ;
        RECT 94.400 21.100 94.800 22.800 ;
        RECT 96.600 21.100 97.000 25.300 ;
        RECT 99.900 25.200 101.100 25.500 ;
        RECT 99.900 23.100 100.200 25.200 ;
        RECT 101.500 25.100 101.800 25.800 ;
        RECT 99.800 21.100 100.200 23.100 ;
        RECT 101.400 21.100 101.800 25.100 ;
        RECT 102.200 27.700 102.600 29.900 ;
        RECT 104.300 29.200 104.900 29.900 ;
        RECT 104.300 28.900 105.000 29.200 ;
        RECT 106.600 28.900 107.000 29.900 ;
        RECT 108.800 29.200 109.200 29.900 ;
        RECT 108.800 28.900 109.800 29.200 ;
        RECT 104.600 28.500 105.000 28.900 ;
        RECT 106.700 28.600 107.000 28.900 ;
        RECT 106.700 28.300 108.100 28.600 ;
        RECT 107.700 28.200 108.100 28.300 ;
        RECT 105.400 27.800 105.800 28.200 ;
        RECT 108.600 27.800 109.000 28.600 ;
        RECT 109.400 28.500 109.800 28.900 ;
        RECT 103.700 27.700 104.100 27.800 ;
        RECT 102.200 27.400 104.100 27.700 ;
        RECT 102.200 25.700 102.600 27.400 ;
        RECT 105.400 27.200 105.700 27.800 ;
        RECT 105.400 27.100 106.100 27.200 ;
        RECT 108.600 27.100 108.900 27.800 ;
        RECT 111.000 27.500 111.400 29.900 ;
        RECT 111.800 27.700 112.200 29.900 ;
        RECT 113.900 29.200 114.500 29.900 ;
        RECT 113.900 28.900 114.600 29.200 ;
        RECT 116.200 28.900 116.600 29.900 ;
        RECT 118.400 29.200 118.800 29.900 ;
        RECT 118.400 28.900 119.400 29.200 ;
        RECT 114.200 28.500 114.600 28.900 ;
        RECT 116.300 28.600 116.600 28.900 ;
        RECT 116.300 28.300 117.700 28.600 ;
        RECT 117.300 28.200 117.700 28.300 ;
        RECT 118.200 27.800 118.600 28.600 ;
        RECT 119.000 28.500 119.400 28.900 ;
        RECT 113.300 27.700 113.700 27.800 ;
        RECT 111.800 27.400 113.700 27.700 ;
        RECT 110.200 27.100 111.000 27.200 ;
        RECT 105.400 26.800 111.000 27.100 ;
        RECT 104.600 26.400 105.000 26.500 ;
        RECT 103.100 26.100 105.000 26.400 ;
        RECT 103.100 26.000 103.500 26.100 ;
        RECT 103.900 25.700 104.300 25.800 ;
        RECT 102.200 25.400 104.300 25.700 ;
        RECT 102.200 21.100 102.600 25.400 ;
        RECT 105.500 25.200 105.800 26.800 ;
        RECT 109.100 26.700 109.500 26.800 ;
        RECT 108.600 26.200 109.000 26.300 ;
        RECT 109.900 26.200 110.300 26.300 ;
        RECT 107.800 25.900 110.300 26.200 ;
        RECT 107.800 25.800 108.200 25.900 ;
        RECT 111.800 25.700 112.200 27.400 ;
        RECT 115.300 27.100 115.700 27.200 ;
        RECT 118.200 27.100 118.500 27.800 ;
        RECT 120.600 27.500 121.000 29.900 ;
        RECT 121.400 27.800 121.800 28.600 ;
        RECT 119.800 27.100 120.600 27.200 ;
        RECT 115.100 26.800 120.600 27.100 ;
        RECT 114.200 26.400 114.600 26.500 ;
        RECT 112.700 26.100 114.600 26.400 ;
        RECT 112.700 26.000 113.100 26.100 ;
        RECT 113.500 25.700 113.900 25.800 ;
        RECT 108.600 25.500 111.400 25.600 ;
        RECT 108.500 25.400 111.400 25.500 ;
        RECT 104.600 24.900 105.800 25.200 ;
        RECT 106.500 25.300 111.400 25.400 ;
        RECT 106.500 25.100 108.900 25.300 ;
        RECT 104.600 24.400 104.900 24.900 ;
        RECT 104.200 24.000 104.900 24.400 ;
        RECT 105.700 24.500 106.100 24.600 ;
        RECT 106.500 24.500 106.800 25.100 ;
        RECT 105.700 24.200 106.800 24.500 ;
        RECT 107.100 24.500 109.800 24.800 ;
        RECT 107.100 24.400 107.500 24.500 ;
        RECT 109.400 24.400 109.800 24.500 ;
        RECT 106.300 23.700 106.700 23.800 ;
        RECT 107.700 23.700 108.100 23.800 ;
        RECT 104.600 23.100 105.000 23.500 ;
        RECT 106.300 23.400 108.100 23.700 ;
        RECT 106.700 23.100 107.000 23.400 ;
        RECT 109.400 23.100 109.800 23.500 ;
        RECT 104.300 21.100 104.900 23.100 ;
        RECT 106.600 21.100 107.000 23.100 ;
        RECT 108.800 22.800 109.800 23.100 ;
        RECT 108.800 21.100 109.200 22.800 ;
        RECT 111.000 21.100 111.400 25.300 ;
        RECT 111.800 25.400 113.900 25.700 ;
        RECT 111.800 21.100 112.200 25.400 ;
        RECT 115.100 25.200 115.400 26.800 ;
        RECT 118.700 26.700 119.100 26.800 ;
        RECT 119.500 26.200 119.900 26.300 ;
        RECT 117.400 25.900 119.900 26.200 ;
        RECT 117.400 25.800 117.800 25.900 ;
        RECT 118.200 25.500 121.000 25.600 ;
        RECT 118.100 25.400 121.000 25.500 ;
        RECT 114.200 24.900 115.400 25.200 ;
        RECT 116.100 25.300 121.000 25.400 ;
        RECT 116.100 25.100 118.500 25.300 ;
        RECT 114.200 24.400 114.500 24.900 ;
        RECT 113.800 24.200 114.500 24.400 ;
        RECT 115.300 24.500 115.700 24.600 ;
        RECT 116.100 24.500 116.400 25.100 ;
        RECT 115.300 24.200 116.400 24.500 ;
        RECT 116.700 24.500 119.400 24.800 ;
        RECT 116.700 24.400 117.100 24.500 ;
        RECT 119.000 24.400 119.400 24.500 ;
        RECT 113.400 24.000 114.500 24.200 ;
        RECT 113.400 23.800 114.100 24.000 ;
        RECT 115.900 23.700 116.300 23.800 ;
        RECT 117.300 23.700 117.700 23.800 ;
        RECT 114.200 23.100 114.600 23.500 ;
        RECT 115.900 23.400 117.700 23.700 ;
        RECT 116.300 23.100 116.600 23.400 ;
        RECT 119.000 23.100 119.400 23.500 ;
        RECT 113.900 21.100 114.500 23.100 ;
        RECT 116.200 21.100 116.600 23.100 ;
        RECT 118.400 22.800 119.400 23.100 ;
        RECT 118.400 21.100 118.800 22.800 ;
        RECT 120.600 21.100 121.000 25.300 ;
        RECT 122.200 21.100 122.600 29.900 ;
        RECT 123.800 27.600 124.200 29.900 ;
        RECT 125.400 27.600 125.800 29.900 ;
        RECT 127.000 27.600 127.400 29.900 ;
        RECT 128.600 27.600 129.000 29.900 ;
        RECT 130.200 27.800 130.600 28.600 ;
        RECT 131.000 28.100 131.400 29.900 ;
        RECT 132.600 28.900 133.000 29.900 ;
        RECT 131.800 28.100 132.200 28.600 ;
        RECT 131.000 27.800 132.200 28.100 ;
        RECT 123.000 27.200 124.200 27.600 ;
        RECT 124.700 27.200 125.800 27.600 ;
        RECT 126.300 27.200 127.400 27.600 ;
        RECT 128.100 27.200 129.000 27.600 ;
        RECT 123.000 25.800 123.400 27.200 ;
        RECT 124.700 26.900 125.100 27.200 ;
        RECT 126.300 26.900 126.700 27.200 ;
        RECT 128.100 26.900 128.500 27.200 ;
        RECT 123.800 26.500 125.100 26.900 ;
        RECT 125.500 26.500 126.700 26.900 ;
        RECT 127.200 26.500 128.500 26.900 ;
        RECT 124.700 25.800 125.100 26.500 ;
        RECT 126.300 25.800 126.700 26.500 ;
        RECT 128.100 25.800 128.500 26.500 ;
        RECT 123.000 25.400 124.200 25.800 ;
        RECT 124.700 25.400 125.800 25.800 ;
        RECT 126.300 25.400 127.400 25.800 ;
        RECT 128.100 25.400 129.000 25.800 ;
        RECT 123.800 21.100 124.200 25.400 ;
        RECT 125.400 21.100 125.800 25.400 ;
        RECT 127.000 21.100 127.400 25.400 ;
        RECT 128.600 21.100 129.000 25.400 ;
        RECT 131.000 21.100 131.400 27.800 ;
        RECT 132.700 27.200 133.000 28.900 ;
        RECT 134.200 27.500 134.600 29.900 ;
        RECT 136.400 29.200 136.800 29.900 ;
        RECT 135.800 28.900 136.800 29.200 ;
        RECT 138.600 28.900 139.000 29.900 ;
        RECT 140.700 29.200 141.300 29.900 ;
        RECT 140.600 28.900 141.300 29.200 ;
        RECT 135.800 28.500 136.200 28.900 ;
        RECT 138.600 28.600 138.900 28.900 ;
        RECT 136.600 28.200 137.000 28.600 ;
        RECT 137.500 28.300 138.900 28.600 ;
        RECT 140.600 28.500 141.000 28.900 ;
        RECT 137.500 28.200 137.900 28.300 ;
        RECT 132.600 26.800 133.000 27.200 ;
        RECT 134.600 27.100 135.400 27.200 ;
        RECT 136.700 27.100 137.000 28.200 ;
        RECT 141.500 27.700 141.900 27.800 ;
        RECT 143.000 27.700 143.400 29.900 ;
        RECT 141.500 27.400 143.400 27.700 ;
        RECT 145.400 27.500 145.800 29.900 ;
        RECT 147.600 29.200 148.000 29.900 ;
        RECT 147.000 28.900 148.000 29.200 ;
        RECT 149.800 28.900 150.200 29.900 ;
        RECT 151.900 29.200 152.500 29.900 ;
        RECT 151.800 28.900 152.500 29.200 ;
        RECT 147.000 28.500 147.400 28.900 ;
        RECT 149.800 28.600 150.100 28.900 ;
        RECT 147.800 28.200 148.200 28.600 ;
        RECT 148.700 28.300 150.100 28.600 ;
        RECT 151.800 28.500 152.200 28.900 ;
        RECT 148.700 28.200 149.100 28.300 ;
        RECT 139.500 27.100 139.900 27.200 ;
        RECT 134.600 26.800 140.100 27.100 ;
        RECT 132.700 25.100 133.000 26.800 ;
        RECT 136.100 26.700 136.500 26.800 ;
        RECT 135.300 26.200 135.700 26.300 ;
        RECT 133.400 25.400 133.800 26.200 ;
        RECT 135.300 25.900 137.800 26.200 ;
        RECT 137.400 25.800 137.800 25.900 ;
        RECT 134.200 25.500 137.000 25.600 ;
        RECT 134.200 25.400 137.100 25.500 ;
        RECT 134.200 25.300 139.100 25.400 ;
        RECT 132.600 24.700 133.500 25.100 ;
        RECT 133.100 21.100 133.500 24.700 ;
        RECT 134.200 21.100 134.600 25.300 ;
        RECT 136.700 25.100 139.100 25.300 ;
        RECT 135.800 24.500 138.500 24.800 ;
        RECT 135.800 24.400 136.200 24.500 ;
        RECT 138.100 24.400 138.500 24.500 ;
        RECT 138.800 24.500 139.100 25.100 ;
        RECT 139.800 25.200 140.100 26.800 ;
        RECT 140.600 26.400 141.000 26.500 ;
        RECT 140.600 26.100 142.500 26.400 ;
        RECT 142.100 26.000 142.500 26.100 ;
        RECT 141.300 25.700 141.700 25.800 ;
        RECT 143.000 25.700 143.400 27.400 ;
        RECT 144.600 27.100 145.000 27.200 ;
        RECT 145.800 27.100 146.600 27.200 ;
        RECT 147.900 27.100 148.200 28.200 ;
        RECT 152.700 27.700 153.100 27.800 ;
        RECT 154.200 27.700 154.600 29.900 ;
        RECT 152.700 27.400 154.600 27.700 ;
        RECT 155.000 27.500 155.400 29.900 ;
        RECT 157.200 29.200 157.600 29.900 ;
        RECT 156.600 28.900 157.600 29.200 ;
        RECT 159.400 28.900 159.800 29.900 ;
        RECT 161.500 29.200 162.100 29.900 ;
        RECT 161.400 28.900 162.100 29.200 ;
        RECT 156.600 28.500 157.000 28.900 ;
        RECT 159.400 28.600 159.700 28.900 ;
        RECT 157.400 28.200 157.800 28.600 ;
        RECT 158.300 28.300 159.700 28.600 ;
        RECT 161.400 28.500 161.800 28.900 ;
        RECT 158.300 28.200 158.700 28.300 ;
        RECT 150.700 27.100 151.100 27.200 ;
        RECT 144.600 26.800 151.300 27.100 ;
        RECT 147.300 26.700 147.700 26.800 ;
        RECT 146.500 26.200 146.900 26.300 ;
        RECT 146.500 25.900 149.000 26.200 ;
        RECT 148.600 25.800 149.000 25.900 ;
        RECT 141.300 25.400 143.400 25.700 ;
        RECT 139.800 24.900 141.000 25.200 ;
        RECT 139.500 24.500 139.900 24.600 ;
        RECT 138.800 24.200 139.900 24.500 ;
        RECT 140.700 24.400 141.000 24.900 ;
        RECT 140.700 24.200 141.400 24.400 ;
        RECT 140.700 24.000 141.800 24.200 ;
        RECT 141.100 23.800 141.800 24.000 ;
        RECT 137.500 23.700 137.900 23.800 ;
        RECT 138.900 23.700 139.300 23.800 ;
        RECT 135.800 23.100 136.200 23.500 ;
        RECT 137.500 23.400 139.300 23.700 ;
        RECT 138.600 23.100 138.900 23.400 ;
        RECT 140.600 23.100 141.000 23.500 ;
        RECT 135.800 22.800 136.800 23.100 ;
        RECT 136.400 21.100 136.800 22.800 ;
        RECT 138.600 21.100 139.000 23.100 ;
        RECT 140.700 21.100 141.300 23.100 ;
        RECT 143.000 21.100 143.400 25.400 ;
        RECT 145.400 25.500 148.200 25.600 ;
        RECT 145.400 25.400 148.300 25.500 ;
        RECT 145.400 25.300 150.300 25.400 ;
        RECT 145.400 21.100 145.800 25.300 ;
        RECT 147.900 25.100 150.300 25.300 ;
        RECT 147.000 24.500 149.700 24.800 ;
        RECT 147.000 24.400 147.400 24.500 ;
        RECT 149.300 24.400 149.700 24.500 ;
        RECT 150.000 24.500 150.300 25.100 ;
        RECT 151.000 25.200 151.300 26.800 ;
        RECT 151.800 26.400 152.200 26.500 ;
        RECT 151.800 26.100 153.700 26.400 ;
        RECT 153.300 26.000 153.700 26.100 ;
        RECT 152.500 25.700 152.900 25.800 ;
        RECT 154.200 25.700 154.600 27.400 ;
        RECT 155.400 27.100 156.200 27.200 ;
        RECT 157.500 27.100 157.800 28.200 ;
        RECT 162.200 27.800 162.600 28.200 ;
        RECT 162.200 27.700 162.700 27.800 ;
        RECT 163.800 27.700 164.200 29.900 ;
        RECT 164.600 27.900 165.000 29.900 ;
        RECT 165.400 28.000 165.800 29.900 ;
        RECT 167.000 28.000 167.400 29.900 ;
        RECT 165.400 27.900 167.400 28.000 ;
        RECT 162.200 27.400 164.200 27.700 ;
        RECT 160.300 27.100 160.700 27.200 ;
        RECT 155.400 26.800 160.900 27.100 ;
        RECT 156.900 26.700 157.300 26.800 ;
        RECT 156.100 26.200 156.500 26.300 ;
        RECT 157.400 26.200 157.800 26.300 ;
        RECT 156.100 25.900 158.600 26.200 ;
        RECT 158.200 25.800 158.600 25.900 ;
        RECT 159.800 26.100 160.200 26.200 ;
        RECT 160.600 26.100 160.900 26.800 ;
        RECT 161.400 26.400 161.800 26.500 ;
        RECT 161.400 26.100 163.300 26.400 ;
        RECT 159.800 25.800 160.900 26.100 ;
        RECT 162.900 26.000 163.300 26.100 ;
        RECT 152.500 25.400 154.600 25.700 ;
        RECT 151.000 24.900 152.200 25.200 ;
        RECT 150.700 24.500 151.100 24.600 ;
        RECT 150.000 24.200 151.100 24.500 ;
        RECT 151.900 24.400 152.200 24.900 ;
        RECT 151.900 24.000 152.600 24.400 ;
        RECT 148.700 23.700 149.100 23.800 ;
        RECT 150.100 23.700 150.500 23.800 ;
        RECT 147.000 23.100 147.400 23.500 ;
        RECT 148.700 23.400 150.500 23.700 ;
        RECT 149.800 23.100 150.100 23.400 ;
        RECT 151.800 23.100 152.200 23.500 ;
        RECT 147.000 22.800 148.000 23.100 ;
        RECT 147.600 21.100 148.000 22.800 ;
        RECT 149.800 21.100 150.200 23.100 ;
        RECT 151.900 21.100 152.500 23.100 ;
        RECT 154.200 21.100 154.600 25.400 ;
        RECT 155.000 25.500 157.800 25.600 ;
        RECT 155.000 25.400 157.900 25.500 ;
        RECT 155.000 25.300 159.900 25.400 ;
        RECT 155.000 21.100 155.400 25.300 ;
        RECT 157.500 25.100 159.900 25.300 ;
        RECT 156.600 24.500 159.300 24.800 ;
        RECT 156.600 24.400 157.000 24.500 ;
        RECT 158.900 24.400 159.300 24.500 ;
        RECT 159.600 24.500 159.900 25.100 ;
        RECT 160.600 25.200 160.900 25.800 ;
        RECT 162.100 25.700 162.500 25.800 ;
        RECT 163.800 25.700 164.200 27.400 ;
        RECT 164.700 27.200 165.000 27.900 ;
        RECT 165.500 27.700 167.300 27.900 ;
        RECT 167.800 27.700 168.200 29.900 ;
        RECT 169.900 29.200 170.500 29.900 ;
        RECT 169.900 28.900 170.600 29.200 ;
        RECT 172.200 28.900 172.600 29.900 ;
        RECT 174.400 29.200 174.800 29.900 ;
        RECT 174.400 28.900 175.400 29.200 ;
        RECT 170.200 28.500 170.600 28.900 ;
        RECT 172.300 28.600 172.600 28.900 ;
        RECT 172.300 28.300 173.700 28.600 ;
        RECT 173.300 28.200 173.700 28.300 ;
        RECT 174.200 28.200 174.600 28.600 ;
        RECT 175.000 28.500 175.400 28.900 ;
        RECT 169.300 27.700 169.700 27.800 ;
        RECT 167.800 27.400 169.700 27.700 ;
        RECT 166.600 27.200 167.000 27.400 ;
        RECT 164.600 26.800 165.900 27.200 ;
        RECT 166.600 26.900 167.400 27.200 ;
        RECT 167.000 26.800 167.400 26.900 ;
        RECT 162.100 25.400 164.200 25.700 ;
        RECT 160.600 24.900 161.800 25.200 ;
        RECT 160.300 24.500 160.700 24.600 ;
        RECT 159.600 24.200 160.700 24.500 ;
        RECT 161.500 24.400 161.800 24.900 ;
        RECT 161.500 24.000 162.200 24.400 ;
        RECT 158.300 23.700 158.700 23.800 ;
        RECT 159.700 23.700 160.100 23.800 ;
        RECT 156.600 23.100 157.000 23.500 ;
        RECT 158.300 23.400 160.100 23.700 ;
        RECT 159.400 23.100 159.700 23.400 ;
        RECT 161.400 23.100 161.800 23.500 ;
        RECT 156.600 22.800 157.600 23.100 ;
        RECT 157.200 21.100 157.600 22.800 ;
        RECT 159.400 21.100 159.800 23.100 ;
        RECT 161.500 21.100 162.100 23.100 ;
        RECT 163.800 21.100 164.200 25.400 ;
        RECT 164.600 25.100 165.000 25.200 ;
        RECT 165.600 25.100 165.900 26.800 ;
        RECT 166.200 26.100 166.600 26.600 ;
        RECT 167.800 26.100 168.200 27.400 ;
        RECT 168.600 26.800 169.000 27.400 ;
        RECT 171.300 27.100 171.700 27.200 ;
        RECT 174.200 27.100 174.500 28.200 ;
        RECT 176.600 27.500 177.000 29.900 ;
        RECT 178.200 28.800 178.600 29.900 ;
        RECT 177.400 27.800 177.800 28.600 ;
        RECT 178.300 27.200 178.600 28.800 ;
        RECT 179.800 27.500 180.200 29.900 ;
        RECT 182.000 29.200 182.400 29.900 ;
        RECT 181.400 28.900 182.400 29.200 ;
        RECT 184.200 28.900 184.600 29.900 ;
        RECT 186.300 29.200 186.900 29.900 ;
        RECT 186.200 28.900 186.900 29.200 ;
        RECT 181.400 28.500 181.800 28.900 ;
        RECT 184.200 28.600 184.500 28.900 ;
        RECT 182.200 28.200 182.600 28.600 ;
        RECT 183.100 28.300 184.500 28.600 ;
        RECT 186.200 28.500 186.600 28.900 ;
        RECT 183.100 28.200 183.500 28.300 ;
        RECT 175.800 27.100 176.600 27.200 ;
        RECT 171.100 26.800 176.600 27.100 ;
        RECT 178.200 26.800 178.600 27.200 ;
        RECT 180.200 27.100 181.000 27.200 ;
        RECT 182.300 27.100 182.600 28.200 ;
        RECT 187.100 27.700 187.500 27.800 ;
        RECT 188.600 27.700 189.000 29.900 ;
        RECT 187.100 27.400 189.000 27.700 ;
        RECT 185.100 27.100 185.500 27.200 ;
        RECT 180.200 26.800 185.700 27.100 ;
        RECT 170.200 26.400 170.600 26.500 ;
        RECT 166.200 25.800 168.200 26.100 ;
        RECT 168.700 26.100 170.600 26.400 ;
        RECT 171.100 26.200 171.400 26.800 ;
        RECT 174.700 26.700 175.100 26.800 ;
        RECT 174.200 26.200 174.600 26.300 ;
        RECT 175.500 26.200 175.900 26.300 ;
        RECT 168.700 26.000 169.100 26.100 ;
        RECT 171.000 25.800 171.400 26.200 ;
        RECT 173.400 25.900 175.900 26.200 ;
        RECT 173.400 25.800 173.800 25.900 ;
        RECT 167.800 25.700 168.200 25.800 ;
        RECT 169.500 25.700 169.900 25.800 ;
        RECT 167.800 25.400 169.900 25.700 ;
        RECT 164.600 24.800 165.300 25.100 ;
        RECT 165.600 24.800 166.100 25.100 ;
        RECT 165.000 24.200 165.300 24.800 ;
        RECT 165.000 23.800 165.400 24.200 ;
        RECT 165.700 21.100 166.100 24.800 ;
        RECT 167.800 21.100 168.200 25.400 ;
        RECT 171.100 25.200 171.400 25.800 ;
        RECT 174.200 25.500 177.000 25.600 ;
        RECT 174.100 25.400 177.000 25.500 ;
        RECT 170.200 24.900 171.400 25.200 ;
        RECT 172.100 25.300 177.000 25.400 ;
        RECT 172.100 25.100 174.500 25.300 ;
        RECT 170.200 24.400 170.500 24.900 ;
        RECT 169.800 24.000 170.500 24.400 ;
        RECT 171.300 24.500 171.700 24.600 ;
        RECT 172.100 24.500 172.400 25.100 ;
        RECT 171.300 24.200 172.400 24.500 ;
        RECT 172.700 24.500 175.400 24.800 ;
        RECT 172.700 24.400 173.100 24.500 ;
        RECT 175.000 24.400 175.400 24.500 ;
        RECT 171.900 23.700 172.300 23.800 ;
        RECT 173.300 23.700 173.700 23.800 ;
        RECT 170.200 23.100 170.600 23.500 ;
        RECT 171.900 23.400 173.700 23.700 ;
        RECT 172.300 23.100 172.600 23.400 ;
        RECT 175.000 23.100 175.400 23.500 ;
        RECT 169.900 21.100 170.500 23.100 ;
        RECT 172.200 21.100 172.600 23.100 ;
        RECT 174.400 22.800 175.400 23.100 ;
        RECT 174.400 21.100 174.800 22.800 ;
        RECT 176.600 21.100 177.000 25.300 ;
        RECT 178.300 25.100 178.600 26.800 ;
        RECT 181.700 26.700 182.100 26.800 ;
        RECT 180.900 26.200 181.300 26.300 ;
        RECT 182.200 26.200 182.600 26.300 ;
        RECT 179.000 25.400 179.400 26.200 ;
        RECT 180.900 25.900 183.400 26.200 ;
        RECT 183.000 25.800 183.400 25.900 ;
        RECT 179.800 25.500 182.600 25.600 ;
        RECT 179.800 25.400 182.700 25.500 ;
        RECT 179.800 25.300 184.700 25.400 ;
        RECT 178.200 24.700 179.100 25.100 ;
        RECT 178.700 21.100 179.100 24.700 ;
        RECT 179.800 21.100 180.200 25.300 ;
        RECT 182.300 25.100 184.700 25.300 ;
        RECT 181.400 24.500 184.100 24.800 ;
        RECT 181.400 24.400 181.800 24.500 ;
        RECT 183.700 24.400 184.100 24.500 ;
        RECT 184.400 24.500 184.700 25.100 ;
        RECT 185.400 25.200 185.700 26.800 ;
        RECT 186.200 26.400 186.600 26.500 ;
        RECT 186.200 26.100 188.100 26.400 ;
        RECT 187.700 26.000 188.100 26.100 ;
        RECT 186.900 25.700 187.300 25.800 ;
        RECT 188.600 25.700 189.000 27.400 ;
        RECT 186.900 25.400 189.000 25.700 ;
        RECT 185.400 24.900 186.600 25.200 ;
        RECT 185.100 24.500 185.500 24.600 ;
        RECT 184.400 24.200 185.500 24.500 ;
        RECT 186.300 24.400 186.600 24.900 ;
        RECT 186.300 24.000 187.000 24.400 ;
        RECT 183.100 23.700 183.500 23.800 ;
        RECT 184.500 23.700 184.900 23.800 ;
        RECT 181.400 23.100 181.800 23.500 ;
        RECT 183.100 23.400 184.900 23.700 ;
        RECT 184.200 23.100 184.500 23.400 ;
        RECT 186.200 23.100 186.600 23.500 ;
        RECT 181.400 22.800 182.400 23.100 ;
        RECT 182.000 21.100 182.400 22.800 ;
        RECT 184.200 21.100 184.600 23.100 ;
        RECT 186.300 21.100 186.900 23.100 ;
        RECT 188.600 21.100 189.000 25.400 ;
        RECT 189.400 26.200 189.800 29.900 ;
        RECT 191.000 27.600 191.400 29.900 ;
        RECT 190.300 27.300 191.400 27.600 ;
        RECT 191.800 27.600 192.200 29.900 ;
        RECT 191.800 27.300 192.900 27.600 ;
        RECT 189.400 25.100 189.700 26.200 ;
        RECT 190.300 25.800 190.600 27.300 ;
        RECT 190.000 25.400 190.600 25.800 ;
        RECT 190.300 25.100 190.600 25.400 ;
        RECT 192.600 25.800 192.900 27.300 ;
        RECT 193.400 26.200 193.800 29.900 ;
        RECT 192.600 25.400 193.200 25.800 ;
        RECT 192.600 25.100 192.900 25.400 ;
        RECT 193.500 25.100 193.800 26.200 ;
        RECT 189.400 21.100 189.800 25.100 ;
        RECT 190.300 24.800 191.400 25.100 ;
        RECT 191.000 21.100 191.400 24.800 ;
        RECT 191.800 24.800 192.900 25.100 ;
        RECT 191.800 21.100 192.200 24.800 ;
        RECT 193.400 21.100 193.800 25.100 ;
        RECT 2.200 16.200 2.600 19.900 ;
        RECT 1.500 15.900 2.600 16.200 ;
        RECT 1.500 15.600 1.800 15.900 ;
        RECT 1.200 15.200 1.800 15.600 ;
        RECT 1.500 13.700 1.800 15.200 ;
        RECT 3.000 15.600 3.400 19.900 ;
        RECT 5.100 17.900 5.700 19.900 ;
        RECT 7.400 17.900 7.800 19.900 ;
        RECT 9.600 18.200 10.000 19.900 ;
        RECT 9.600 17.900 10.600 18.200 ;
        RECT 5.400 17.500 5.800 17.900 ;
        RECT 7.500 17.600 7.800 17.900 ;
        RECT 7.100 17.300 8.900 17.600 ;
        RECT 10.200 17.500 10.600 17.900 ;
        RECT 7.100 17.200 7.500 17.300 ;
        RECT 8.500 17.200 8.900 17.300 ;
        RECT 5.000 16.600 5.700 17.000 ;
        RECT 5.400 16.100 5.700 16.600 ;
        RECT 6.500 16.500 7.600 16.800 ;
        RECT 6.500 16.400 6.900 16.500 ;
        RECT 5.400 15.800 6.600 16.100 ;
        RECT 3.000 15.300 5.100 15.600 ;
        RECT 1.500 13.400 2.600 13.700 ;
        RECT 2.200 11.100 2.600 13.400 ;
        RECT 3.000 13.600 3.400 15.300 ;
        RECT 4.700 15.200 5.100 15.300 ;
        RECT 3.900 14.900 4.300 15.000 ;
        RECT 3.900 14.600 5.800 14.900 ;
        RECT 5.400 14.500 5.800 14.600 ;
        RECT 6.300 14.200 6.600 15.800 ;
        RECT 7.300 15.900 7.600 16.500 ;
        RECT 7.900 16.500 8.300 16.600 ;
        RECT 10.200 16.500 10.600 16.600 ;
        RECT 7.900 16.200 10.600 16.500 ;
        RECT 7.300 15.700 9.700 15.900 ;
        RECT 11.800 15.700 12.200 19.900 ;
        RECT 12.900 16.300 13.300 19.900 ;
        RECT 12.900 15.900 13.800 16.300 ;
        RECT 7.300 15.600 12.200 15.700 ;
        RECT 9.300 15.500 12.200 15.600 ;
        RECT 9.400 15.400 12.200 15.500 ;
        RECT 8.600 15.100 9.000 15.200 ;
        RECT 8.600 14.800 11.100 15.100 ;
        RECT 12.600 14.800 13.000 15.600 ;
        RECT 10.700 14.700 11.100 14.800 ;
        RECT 9.900 14.200 10.300 14.300 ;
        RECT 13.400 14.200 13.700 15.900 ;
        RECT 15.000 15.700 15.400 19.900 ;
        RECT 17.200 18.200 17.600 19.900 ;
        RECT 16.600 17.900 17.600 18.200 ;
        RECT 19.400 17.900 19.800 19.900 ;
        RECT 21.500 17.900 22.100 19.900 ;
        RECT 16.600 17.500 17.000 17.900 ;
        RECT 19.400 17.600 19.700 17.900 ;
        RECT 18.300 17.300 20.100 17.600 ;
        RECT 21.400 17.500 21.800 17.900 ;
        RECT 18.300 17.200 18.700 17.300 ;
        RECT 19.700 17.200 20.100 17.300 ;
        RECT 16.600 16.500 17.000 16.600 ;
        RECT 18.900 16.500 19.300 16.600 ;
        RECT 16.600 16.200 19.300 16.500 ;
        RECT 19.600 16.500 20.700 16.800 ;
        RECT 19.600 15.900 19.900 16.500 ;
        RECT 20.300 16.400 20.700 16.500 ;
        RECT 21.500 16.600 22.200 17.000 ;
        RECT 21.500 16.100 21.800 16.600 ;
        RECT 17.500 15.700 19.900 15.900 ;
        RECT 15.000 15.600 19.900 15.700 ;
        RECT 20.600 15.800 21.800 16.100 ;
        RECT 15.000 15.500 17.900 15.600 ;
        RECT 15.000 15.400 17.800 15.500 ;
        RECT 20.600 15.200 20.900 15.800 ;
        RECT 23.800 15.600 24.200 19.900 ;
        RECT 24.900 19.200 25.300 19.900 ;
        RECT 24.900 18.800 25.800 19.200 ;
        RECT 24.900 16.300 25.300 18.800 ;
        RECT 24.900 15.900 25.800 16.300 ;
        RECT 27.000 16.200 27.400 19.900 ;
        RECT 28.600 16.200 29.000 19.900 ;
        RECT 27.000 15.900 29.000 16.200 ;
        RECT 29.400 15.900 29.800 19.900 ;
        RECT 22.100 15.300 24.200 15.600 ;
        RECT 22.100 15.200 22.500 15.300 ;
        RECT 18.200 15.100 18.600 15.200 ;
        RECT 16.100 14.800 18.600 15.100 ;
        RECT 20.600 14.800 21.000 15.200 ;
        RECT 22.900 14.900 23.300 15.000 ;
        RECT 16.100 14.700 16.500 14.800 ;
        RECT 17.400 14.700 17.800 14.800 ;
        RECT 16.900 14.200 17.300 14.300 ;
        RECT 20.600 14.200 20.900 14.800 ;
        RECT 21.400 14.600 23.300 14.900 ;
        RECT 21.400 14.500 21.800 14.600 ;
        RECT 6.300 13.900 11.800 14.200 ;
        RECT 6.500 13.800 6.900 13.900 ;
        RECT 3.000 13.300 4.900 13.600 ;
        RECT 3.000 11.100 3.400 13.300 ;
        RECT 4.500 13.200 4.900 13.300 ;
        RECT 9.400 12.800 9.700 13.900 ;
        RECT 11.000 13.800 11.800 13.900 ;
        RECT 13.400 13.800 13.800 14.200 ;
        RECT 15.400 13.900 20.900 14.200 ;
        RECT 15.400 13.800 16.200 13.900 ;
        RECT 8.500 12.700 8.900 12.800 ;
        RECT 5.400 12.100 5.800 12.500 ;
        RECT 7.500 12.400 8.900 12.700 ;
        RECT 9.400 12.400 9.800 12.800 ;
        RECT 7.500 12.100 7.800 12.400 ;
        RECT 10.200 12.100 10.600 12.500 ;
        RECT 5.100 11.800 5.800 12.100 ;
        RECT 5.100 11.100 5.700 11.800 ;
        RECT 7.400 11.100 7.800 12.100 ;
        RECT 9.600 11.800 10.600 12.100 ;
        RECT 9.600 11.100 10.000 11.800 ;
        RECT 11.800 11.100 12.200 13.500 ;
        RECT 13.400 12.200 13.700 13.800 ;
        RECT 14.200 12.400 14.600 13.200 ;
        RECT 13.400 11.100 13.800 12.200 ;
        RECT 15.000 11.100 15.400 13.500 ;
        RECT 17.500 12.800 17.800 13.900 ;
        RECT 20.300 13.800 20.700 13.900 ;
        RECT 23.800 13.600 24.200 15.300 ;
        RECT 24.600 14.800 25.000 15.600 ;
        RECT 22.300 13.300 24.200 13.600 ;
        RECT 22.300 13.200 22.700 13.300 ;
        RECT 16.600 12.100 17.000 12.500 ;
        RECT 17.400 12.400 17.800 12.800 ;
        RECT 18.300 12.700 18.700 12.800 ;
        RECT 18.300 12.400 19.700 12.700 ;
        RECT 19.400 12.100 19.700 12.400 ;
        RECT 21.400 12.100 21.800 12.500 ;
        RECT 16.600 11.800 17.600 12.100 ;
        RECT 17.200 11.100 17.600 11.800 ;
        RECT 19.400 11.100 19.800 12.100 ;
        RECT 21.400 11.800 22.100 12.100 ;
        RECT 21.500 11.100 22.100 11.800 ;
        RECT 23.800 11.100 24.200 13.300 ;
        RECT 25.400 14.200 25.700 15.900 ;
        RECT 27.400 15.200 27.800 15.400 ;
        RECT 29.400 15.200 29.700 15.900 ;
        RECT 27.000 14.900 27.800 15.200 ;
        RECT 28.600 14.900 29.800 15.200 ;
        RECT 27.000 14.800 27.400 14.900 ;
        RECT 25.400 13.800 25.800 14.200 ;
        RECT 27.800 13.800 28.200 14.600 ;
        RECT 25.400 12.100 25.700 13.800 ;
        RECT 28.600 13.200 28.900 14.900 ;
        RECT 29.400 14.800 29.800 14.900 ;
        RECT 30.200 13.400 30.600 14.200 ;
        RECT 26.200 12.400 26.600 13.200 ;
        RECT 25.400 11.100 25.800 12.100 ;
        RECT 28.600 11.100 29.000 13.200 ;
        RECT 29.400 12.800 29.800 13.200 ;
        RECT 31.000 13.100 31.400 19.900 ;
        RECT 31.800 15.800 32.200 16.600 ;
        RECT 33.900 16.300 34.300 19.900 ;
        RECT 33.400 15.900 34.300 16.300 ;
        RECT 33.500 14.200 33.800 15.900 ;
        RECT 35.000 15.600 35.400 19.900 ;
        RECT 37.100 17.900 37.700 19.900 ;
        RECT 39.400 17.900 39.800 19.900 ;
        RECT 41.600 18.200 42.000 19.900 ;
        RECT 41.600 17.900 42.600 18.200 ;
        RECT 37.400 17.500 37.800 17.900 ;
        RECT 39.500 17.600 39.800 17.900 ;
        RECT 39.100 17.300 40.900 17.600 ;
        RECT 42.200 17.500 42.600 17.900 ;
        RECT 39.100 17.200 39.500 17.300 ;
        RECT 40.500 17.200 40.900 17.300 ;
        RECT 36.600 17.000 37.300 17.200 ;
        RECT 36.600 16.800 37.700 17.000 ;
        RECT 37.000 16.600 37.700 16.800 ;
        RECT 37.400 16.100 37.700 16.600 ;
        RECT 38.500 16.500 39.600 16.800 ;
        RECT 38.500 16.400 38.900 16.500 ;
        RECT 37.400 15.800 38.600 16.100 ;
        RECT 34.200 14.800 34.600 15.600 ;
        RECT 35.000 15.300 37.100 15.600 ;
        RECT 33.400 13.800 33.800 14.200 ;
        RECT 32.600 13.100 33.000 13.200 ;
        RECT 33.500 13.100 33.800 13.800 ;
        RECT 35.000 13.600 35.400 15.300 ;
        RECT 36.700 15.200 37.100 15.300 ;
        RECT 35.900 14.900 36.300 15.000 ;
        RECT 35.900 14.600 37.800 14.900 ;
        RECT 37.400 14.500 37.800 14.600 ;
        RECT 38.300 14.200 38.600 15.800 ;
        RECT 39.300 15.900 39.600 16.500 ;
        RECT 39.900 16.500 40.300 16.600 ;
        RECT 42.200 16.500 42.600 16.600 ;
        RECT 39.900 16.200 42.600 16.500 ;
        RECT 39.300 15.700 41.700 15.900 ;
        RECT 43.800 15.700 44.200 19.900 ;
        RECT 47.000 17.900 47.400 19.900 ;
        RECT 39.300 15.600 44.200 15.700 ;
        RECT 41.300 15.500 44.200 15.600 ;
        RECT 47.100 15.800 47.400 17.900 ;
        RECT 48.600 15.900 49.000 19.900 ;
        RECT 47.100 15.500 48.300 15.800 ;
        RECT 41.400 15.400 44.200 15.500 ;
        RECT 40.600 15.100 41.000 15.200 ;
        RECT 40.600 14.800 43.100 15.100 ;
        RECT 47.000 14.800 47.400 15.200 ;
        RECT 42.700 14.700 43.100 14.800 ;
        RECT 41.900 14.200 42.300 14.300 ;
        RECT 38.300 13.900 43.800 14.200 ;
        RECT 38.500 13.800 38.900 13.900 ;
        RECT 35.000 13.300 36.900 13.600 ;
        RECT 34.200 13.100 34.600 13.200 ;
        RECT 31.000 12.800 33.000 13.100 ;
        RECT 33.400 12.800 34.600 13.100 ;
        RECT 29.300 12.400 29.700 12.800 ;
        RECT 31.500 11.100 31.900 12.800 ;
        RECT 32.600 12.400 33.000 12.800 ;
        RECT 33.500 12.100 33.800 12.800 ;
        RECT 33.400 11.100 33.800 12.100 ;
        RECT 35.000 11.100 35.400 13.300 ;
        RECT 36.500 13.200 36.900 13.300 ;
        RECT 41.400 12.800 41.700 13.900 ;
        RECT 43.000 13.800 43.800 13.900 ;
        RECT 46.200 13.800 46.600 14.600 ;
        RECT 47.100 14.400 47.400 14.800 ;
        RECT 47.100 14.100 47.600 14.400 ;
        RECT 47.200 14.000 47.600 14.100 ;
        RECT 48.000 13.800 48.300 15.500 ;
        RECT 48.700 15.200 49.000 15.900 ;
        RECT 48.600 14.800 49.000 15.200 ;
        RECT 48.000 13.700 48.400 13.800 ;
        RECT 46.900 13.500 48.400 13.700 ;
        RECT 40.500 12.700 40.900 12.800 ;
        RECT 37.400 12.100 37.800 12.500 ;
        RECT 39.500 12.400 40.900 12.700 ;
        RECT 41.400 12.400 41.800 12.800 ;
        RECT 39.500 12.100 39.800 12.400 ;
        RECT 42.200 12.100 42.600 12.500 ;
        RECT 37.100 11.800 37.800 12.100 ;
        RECT 37.100 11.100 37.700 11.800 ;
        RECT 39.400 11.100 39.800 12.100 ;
        RECT 41.600 11.800 42.600 12.100 ;
        RECT 41.600 11.100 42.000 11.800 ;
        RECT 43.800 11.100 44.200 13.500 ;
        RECT 46.300 13.400 48.400 13.500 ;
        RECT 46.300 13.200 47.200 13.400 ;
        RECT 46.300 13.100 46.600 13.200 ;
        RECT 48.700 13.100 49.000 14.800 ;
        RECT 46.200 11.100 46.600 13.100 ;
        RECT 48.300 12.600 49.000 13.100 ;
        RECT 49.400 15.600 49.800 19.900 ;
        RECT 51.500 17.900 52.100 19.900 ;
        RECT 53.800 17.900 54.200 19.900 ;
        RECT 56.000 18.200 56.400 19.900 ;
        RECT 56.000 17.900 57.000 18.200 ;
        RECT 51.800 17.500 52.200 17.900 ;
        RECT 53.900 17.600 54.200 17.900 ;
        RECT 53.500 17.300 55.300 17.600 ;
        RECT 56.600 17.500 57.000 17.900 ;
        RECT 53.500 17.200 53.900 17.300 ;
        RECT 54.900 17.200 55.300 17.300 ;
        RECT 51.400 16.600 52.100 17.000 ;
        RECT 51.800 16.100 52.100 16.600 ;
        RECT 52.900 16.500 54.000 16.800 ;
        RECT 52.900 16.400 53.300 16.500 ;
        RECT 51.800 15.800 53.000 16.100 ;
        RECT 49.400 15.300 51.500 15.600 ;
        RECT 49.400 13.600 49.800 15.300 ;
        RECT 51.100 15.200 51.500 15.300 ;
        RECT 50.300 14.900 50.700 15.000 ;
        RECT 50.300 14.600 52.200 14.900 ;
        RECT 51.800 14.500 52.200 14.600 ;
        RECT 52.700 14.200 53.000 15.800 ;
        RECT 53.700 15.900 54.000 16.500 ;
        RECT 54.300 16.500 54.700 16.600 ;
        RECT 56.600 16.500 57.000 16.600 ;
        RECT 54.300 16.200 57.000 16.500 ;
        RECT 53.700 15.700 56.100 15.900 ;
        RECT 58.200 15.700 58.600 19.900 ;
        RECT 53.700 15.600 58.600 15.700 ;
        RECT 59.800 15.600 60.200 19.900 ;
        RECT 61.400 15.600 61.800 19.900 ;
        RECT 63.000 15.600 63.400 19.900 ;
        RECT 64.600 15.600 65.000 19.900 ;
        RECT 55.700 15.500 58.600 15.600 ;
        RECT 55.800 15.400 58.600 15.500 ;
        RECT 59.000 15.200 60.200 15.600 ;
        RECT 60.700 15.200 61.800 15.600 ;
        RECT 62.300 15.200 63.400 15.600 ;
        RECT 64.100 15.200 65.000 15.600 ;
        RECT 66.200 15.700 66.600 19.900 ;
        RECT 68.400 18.200 68.800 19.900 ;
        RECT 67.800 17.900 68.800 18.200 ;
        RECT 70.600 17.900 71.000 19.900 ;
        RECT 72.700 17.900 73.300 19.900 ;
        RECT 67.800 17.500 68.200 17.900 ;
        RECT 70.600 17.600 70.900 17.900 ;
        RECT 69.500 17.300 71.300 17.600 ;
        RECT 72.600 17.500 73.000 17.900 ;
        RECT 69.500 17.200 69.900 17.300 ;
        RECT 70.900 17.200 71.300 17.300 ;
        RECT 67.800 16.500 68.200 16.600 ;
        RECT 70.100 16.500 70.500 16.600 ;
        RECT 67.800 16.200 70.500 16.500 ;
        RECT 70.800 16.500 71.900 16.800 ;
        RECT 70.800 15.900 71.100 16.500 ;
        RECT 71.500 16.400 71.900 16.500 ;
        RECT 72.700 16.600 73.400 17.000 ;
        RECT 72.700 16.100 73.000 16.600 ;
        RECT 68.700 15.700 71.100 15.900 ;
        RECT 66.200 15.600 71.100 15.700 ;
        RECT 71.800 15.800 73.000 16.100 ;
        RECT 66.200 15.500 69.100 15.600 ;
        RECT 66.200 15.400 69.000 15.500 ;
        RECT 55.000 15.100 55.400 15.200 ;
        RECT 55.000 14.800 57.500 15.100 ;
        RECT 57.100 14.700 57.500 14.800 ;
        RECT 56.300 14.200 56.700 14.300 ;
        RECT 52.700 13.900 58.200 14.200 ;
        RECT 52.900 13.800 53.300 13.900 ;
        RECT 49.400 13.300 51.300 13.600 ;
        RECT 48.300 12.200 48.700 12.600 ;
        RECT 48.300 11.800 49.000 12.200 ;
        RECT 48.300 11.100 48.700 11.800 ;
        RECT 49.400 11.100 49.800 13.300 ;
        RECT 50.900 13.200 51.300 13.300 ;
        RECT 55.800 12.800 56.100 13.900 ;
        RECT 57.400 13.800 58.200 13.900 ;
        RECT 59.000 13.800 59.400 15.200 ;
        RECT 60.700 14.500 61.100 15.200 ;
        RECT 62.300 14.500 62.700 15.200 ;
        RECT 64.100 14.500 64.500 15.200 ;
        RECT 69.400 15.100 69.800 15.200 ;
        RECT 67.300 14.800 69.800 15.100 ;
        RECT 67.300 14.700 67.700 14.800 ;
        RECT 59.800 14.100 61.100 14.500 ;
        RECT 61.500 14.100 62.700 14.500 ;
        RECT 63.200 14.100 64.500 14.500 ;
        RECT 68.100 14.200 68.500 14.300 ;
        RECT 71.800 14.200 72.100 15.800 ;
        RECT 75.000 15.600 75.400 19.900 ;
        RECT 73.300 15.300 75.400 15.600 ;
        RECT 73.300 15.200 73.700 15.300 ;
        RECT 74.100 14.900 74.500 15.000 ;
        RECT 72.600 14.600 74.500 14.900 ;
        RECT 72.600 14.500 73.000 14.600 ;
        RECT 60.700 13.800 61.100 14.100 ;
        RECT 62.300 13.800 62.700 14.100 ;
        RECT 64.100 13.800 64.500 14.100 ;
        RECT 66.600 13.900 72.100 14.200 ;
        RECT 66.600 13.800 67.400 13.900 ;
        RECT 54.900 12.700 55.300 12.800 ;
        RECT 51.800 12.100 52.200 12.500 ;
        RECT 53.900 12.400 55.300 12.700 ;
        RECT 55.800 12.400 56.200 12.800 ;
        RECT 53.900 12.100 54.200 12.400 ;
        RECT 56.600 12.100 57.000 12.500 ;
        RECT 51.500 11.800 52.200 12.100 ;
        RECT 51.500 11.100 52.100 11.800 ;
        RECT 53.800 11.100 54.200 12.100 ;
        RECT 56.000 11.800 57.000 12.100 ;
        RECT 56.000 11.100 56.400 11.800 ;
        RECT 58.200 11.100 58.600 13.500 ;
        RECT 59.000 13.400 60.200 13.800 ;
        RECT 60.700 13.400 61.800 13.800 ;
        RECT 62.300 13.400 63.400 13.800 ;
        RECT 64.100 13.400 65.000 13.800 ;
        RECT 59.800 11.100 60.200 13.400 ;
        RECT 61.400 11.100 61.800 13.400 ;
        RECT 63.000 11.100 63.400 13.400 ;
        RECT 64.600 11.100 65.000 13.400 ;
        RECT 66.200 11.100 66.600 13.500 ;
        RECT 68.700 12.800 69.000 13.900 ;
        RECT 71.500 13.800 71.900 13.900 ;
        RECT 75.000 13.600 75.400 15.300 ;
        RECT 73.500 13.300 75.400 13.600 ;
        RECT 73.500 13.200 73.900 13.300 ;
        RECT 67.800 12.100 68.200 12.500 ;
        RECT 68.600 12.400 69.000 12.800 ;
        RECT 69.500 12.700 69.900 12.800 ;
        RECT 69.500 12.400 70.900 12.700 ;
        RECT 70.600 12.100 70.900 12.400 ;
        RECT 72.600 12.100 73.000 12.500 ;
        RECT 67.800 11.800 68.800 12.100 ;
        RECT 68.400 11.100 68.800 11.800 ;
        RECT 70.600 11.100 71.000 12.100 ;
        RECT 72.600 11.800 73.300 12.100 ;
        RECT 72.700 11.100 73.300 11.800 ;
        RECT 75.000 11.100 75.400 13.300 ;
        RECT 75.800 15.900 76.200 19.900 ;
        RECT 77.400 17.900 77.800 19.900 ;
        RECT 75.800 15.200 76.100 15.900 ;
        RECT 77.400 15.800 77.700 17.900 ;
        RECT 78.200 16.100 78.600 16.200 ;
        RECT 79.000 16.100 79.400 16.600 ;
        RECT 78.200 15.800 79.400 16.100 ;
        RECT 76.500 15.500 77.700 15.800 ;
        RECT 75.800 14.800 76.200 15.200 ;
        RECT 75.800 13.100 76.100 14.800 ;
        RECT 76.500 13.800 76.800 15.500 ;
        RECT 77.400 14.800 77.800 15.200 ;
        RECT 77.400 14.400 77.700 14.800 ;
        RECT 77.200 14.100 77.700 14.400 ;
        RECT 78.200 14.100 78.600 14.600 ;
        RECT 79.000 14.100 79.400 14.200 ;
        RECT 77.200 14.000 77.600 14.100 ;
        RECT 78.200 13.800 79.400 14.100 ;
        RECT 76.400 13.700 76.800 13.800 ;
        RECT 76.400 13.500 77.900 13.700 ;
        RECT 76.400 13.400 78.500 13.500 ;
        RECT 77.600 13.200 78.500 13.400 ;
        RECT 78.200 13.100 78.500 13.200 ;
        RECT 79.800 13.100 80.200 19.900 ;
        RECT 81.700 19.200 82.100 19.900 ;
        RECT 81.400 18.800 82.100 19.200 ;
        RECT 81.700 16.300 82.100 18.800 ;
        RECT 81.700 15.900 82.600 16.300 ;
        RECT 81.400 14.800 81.800 15.600 ;
        RECT 82.200 14.200 82.500 15.900 ;
        RECT 84.600 15.100 85.000 19.900 ;
        RECT 85.400 16.200 85.800 19.900 ;
        RECT 87.000 16.200 87.400 19.900 ;
        RECT 85.400 15.900 87.400 16.200 ;
        RECT 87.800 15.900 88.200 19.900 ;
        RECT 89.000 16.800 89.400 17.200 ;
        RECT 89.000 16.200 89.300 16.800 ;
        RECT 89.700 16.200 90.100 19.900 ;
        RECT 92.100 19.200 92.500 19.900 ;
        RECT 91.800 18.800 92.500 19.200 ;
        RECT 88.600 15.900 89.300 16.200 ;
        RECT 89.600 15.900 90.100 16.200 ;
        RECT 92.100 16.300 92.500 18.800 ;
        RECT 92.100 15.900 93.000 16.300 ;
        RECT 94.200 16.200 94.600 19.900 ;
        RECT 94.200 15.900 95.300 16.200 ;
        RECT 95.800 15.900 96.200 19.900 ;
        RECT 98.200 16.900 98.600 19.900 ;
        RECT 98.300 16.600 98.600 16.900 ;
        RECT 99.800 19.600 101.800 19.900 ;
        RECT 99.800 16.900 100.200 19.600 ;
        RECT 100.600 16.900 101.000 19.300 ;
        RECT 101.400 17.000 101.800 19.600 ;
        RECT 102.300 19.600 104.100 19.900 ;
        RECT 102.300 19.500 102.600 19.600 ;
        RECT 99.800 16.600 100.100 16.900 ;
        RECT 98.300 16.300 100.100 16.600 ;
        RECT 100.700 16.700 101.000 16.900 ;
        RECT 102.200 16.700 102.600 19.500 ;
        RECT 103.800 19.500 104.100 19.600 ;
        RECT 100.700 16.500 102.600 16.700 ;
        RECT 103.000 16.500 103.400 19.300 ;
        RECT 103.800 16.500 104.200 19.500 ;
        RECT 100.700 16.400 102.500 16.500 ;
        RECT 103.000 16.200 103.300 16.500 ;
        RECT 103.000 16.100 103.400 16.200 ;
        RECT 85.800 15.200 86.200 15.400 ;
        RECT 87.800 15.200 88.100 15.900 ;
        RECT 88.600 15.800 89.000 15.900 ;
        RECT 85.400 15.100 86.200 15.200 ;
        RECT 84.600 14.900 86.200 15.100 ;
        RECT 87.000 14.900 88.200 15.200 ;
        RECT 84.600 14.800 85.800 14.900 ;
        RECT 80.600 13.400 81.000 14.200 ;
        RECT 82.200 13.800 82.600 14.200 ;
        RECT 75.800 12.600 76.500 13.100 ;
        RECT 76.100 11.100 76.500 12.600 ;
        RECT 78.200 11.100 78.600 13.100 ;
        RECT 79.300 12.800 80.200 13.100 ;
        RECT 79.300 11.100 79.700 12.800 ;
        RECT 82.200 12.100 82.500 13.800 ;
        RECT 83.000 12.400 83.400 13.200 ;
        RECT 83.800 12.400 84.200 13.200 ;
        RECT 82.200 11.100 82.600 12.100 ;
        RECT 84.600 11.100 85.000 14.800 ;
        RECT 86.200 13.800 86.600 14.600 ;
        RECT 87.000 13.100 87.300 14.900 ;
        RECT 87.800 14.800 88.200 14.900 ;
        RECT 89.600 14.200 89.900 15.900 ;
        RECT 90.200 14.400 90.600 15.200 ;
        RECT 91.800 14.800 92.200 15.600 ;
        RECT 92.600 14.200 92.900 15.900 ;
        RECT 95.000 15.600 95.300 15.900 ;
        RECT 95.000 15.200 95.600 15.600 ;
        RECT 88.600 13.800 89.900 14.200 ;
        RECT 91.000 14.100 91.400 14.200 ;
        RECT 90.600 13.800 91.400 14.100 ;
        RECT 92.600 13.800 93.000 14.200 ;
        RECT 87.800 13.100 88.200 13.200 ;
        RECT 88.700 13.100 89.000 13.800 ;
        RECT 90.600 13.600 91.000 13.800 ;
        RECT 89.500 13.100 91.300 13.300 ;
        RECT 87.000 11.100 87.400 13.100 ;
        RECT 87.800 12.800 89.000 13.100 ;
        RECT 87.700 12.400 88.100 12.800 ;
        RECT 88.600 11.100 89.000 12.800 ;
        RECT 89.400 13.000 91.400 13.100 ;
        RECT 89.400 11.100 89.800 13.000 ;
        RECT 91.000 11.100 91.400 13.000 ;
        RECT 92.600 12.100 92.900 13.800 ;
        RECT 95.000 13.700 95.300 15.200 ;
        RECT 95.900 14.800 96.200 15.900 ;
        RECT 101.700 15.800 103.400 16.100 ;
        RECT 100.600 14.800 101.400 15.200 ;
        RECT 94.200 13.400 95.300 13.700 ;
        RECT 93.400 12.400 93.800 13.200 ;
        RECT 92.600 11.100 93.000 12.100 ;
        RECT 94.200 11.100 94.600 13.400 ;
        RECT 95.800 11.100 96.200 14.800 ;
        RECT 99.000 14.100 99.400 14.200 ;
        RECT 99.800 14.100 100.600 14.200 ;
        RECT 99.000 13.800 100.600 14.100 ;
        RECT 99.000 13.100 99.900 13.200 ;
        RECT 100.600 13.100 101.000 13.200 ;
        RECT 99.000 12.800 101.000 13.100 ;
        RECT 101.700 12.500 102.000 15.800 ;
        RECT 105.400 15.100 105.800 19.900 ;
        RECT 106.200 15.800 106.600 16.600 ;
        RECT 108.300 16.200 108.700 19.900 ;
        RECT 111.500 19.200 111.900 19.900 ;
        RECT 111.000 18.800 111.900 19.200 ;
        RECT 109.000 16.800 109.400 17.200 ;
        RECT 109.100 16.200 109.400 16.800 ;
        RECT 111.500 16.300 111.900 18.800 ;
        RECT 108.300 15.900 108.800 16.200 ;
        RECT 109.100 15.900 109.800 16.200 ;
        RECT 111.000 15.900 111.900 16.300 ;
        RECT 112.600 15.900 113.000 19.900 ;
        RECT 113.400 16.200 113.800 19.900 ;
        RECT 115.000 16.200 115.400 19.900 ;
        RECT 113.400 15.900 115.400 16.200 ;
        RECT 107.800 15.100 108.200 15.200 ;
        RECT 105.400 14.800 108.200 15.100 ;
        RECT 103.800 14.100 104.200 14.200 ;
        RECT 104.600 14.100 105.000 14.200 ;
        RECT 103.800 13.800 105.000 14.100 ;
        RECT 104.600 13.400 105.000 13.800 ;
        RECT 105.400 13.100 105.800 14.800 ;
        RECT 107.800 14.400 108.200 14.800 ;
        RECT 108.500 14.200 108.800 15.900 ;
        RECT 109.400 15.800 109.800 15.900 ;
        RECT 111.100 14.200 111.400 15.900 ;
        RECT 111.800 15.100 112.200 15.600 ;
        RECT 112.700 15.200 113.000 15.900 ;
        RECT 114.600 15.200 115.000 15.400 ;
        RECT 112.600 15.100 113.800 15.200 ;
        RECT 111.800 14.900 113.800 15.100 ;
        RECT 114.600 14.900 115.400 15.200 ;
        RECT 111.800 14.800 113.000 14.900 ;
        RECT 107.000 14.100 107.400 14.200 ;
        RECT 107.000 13.800 107.800 14.100 ;
        RECT 108.500 13.800 109.800 14.200 ;
        RECT 111.000 13.800 111.400 14.200 ;
        RECT 107.400 13.600 107.800 13.800 ;
        RECT 107.100 13.100 108.900 13.300 ;
        RECT 109.400 13.100 109.700 13.800 ;
        RECT 110.200 13.100 110.600 13.200 ;
        RECT 105.400 12.800 106.300 13.100 ;
        RECT 100.000 12.200 102.000 12.500 ;
        RECT 105.900 12.200 106.300 12.800 ;
        RECT 99.800 11.800 100.300 12.200 ;
        RECT 101.400 12.100 102.000 12.200 ;
        RECT 99.800 11.100 100.200 11.800 ;
        RECT 101.400 11.100 101.800 12.100 ;
        RECT 105.400 11.800 106.300 12.200 ;
        RECT 105.900 11.100 106.300 11.800 ;
        RECT 107.000 13.000 109.000 13.100 ;
        RECT 107.000 11.100 107.400 13.000 ;
        RECT 108.600 11.100 109.000 13.000 ;
        RECT 109.400 12.800 110.600 13.100 ;
        RECT 109.400 11.100 109.800 12.800 ;
        RECT 110.200 12.400 110.600 12.800 ;
        RECT 111.100 12.100 111.400 13.800 ;
        RECT 111.800 13.100 112.200 13.200 ;
        RECT 112.600 13.100 113.000 13.200 ;
        RECT 113.500 13.100 113.800 14.900 ;
        RECT 115.000 14.800 115.400 14.900 ;
        RECT 114.200 14.100 114.600 14.600 ;
        RECT 115.800 14.100 116.200 19.900 ;
        RECT 117.700 16.300 118.100 19.900 ;
        RECT 117.700 15.900 118.600 16.300 ;
        RECT 117.400 14.800 117.800 15.600 ;
        RECT 114.200 13.800 116.200 14.100 ;
        RECT 111.800 12.800 113.000 13.100 ;
        RECT 112.700 12.400 113.100 12.800 ;
        RECT 111.000 11.100 111.400 12.100 ;
        RECT 113.400 11.100 113.800 13.100 ;
        RECT 115.800 11.100 116.200 13.800 ;
        RECT 116.600 14.100 117.000 14.200 ;
        RECT 117.400 14.100 117.700 14.800 ;
        RECT 116.600 13.800 117.700 14.100 ;
        RECT 118.200 14.200 118.500 15.900 ;
        RECT 119.000 14.800 119.400 15.200 ;
        RECT 118.200 14.100 118.600 14.200 ;
        RECT 119.000 14.100 119.300 14.800 ;
        RECT 118.200 13.800 119.300 14.100 ;
        RECT 116.600 13.400 117.000 13.800 ;
        RECT 118.200 12.100 118.500 13.800 ;
        RECT 119.000 13.100 119.400 13.200 ;
        RECT 119.800 13.100 120.200 19.900 ;
        RECT 121.400 15.600 121.800 19.900 ;
        RECT 123.500 17.900 124.100 19.900 ;
        RECT 125.800 17.900 126.200 19.900 ;
        RECT 128.000 18.200 128.400 19.900 ;
        RECT 128.000 17.900 129.000 18.200 ;
        RECT 123.800 17.500 124.200 17.900 ;
        RECT 125.900 17.600 126.200 17.900 ;
        RECT 125.500 17.300 127.300 17.600 ;
        RECT 128.600 17.500 129.000 17.900 ;
        RECT 125.500 17.200 125.900 17.300 ;
        RECT 126.900 17.200 127.300 17.300 ;
        RECT 123.400 16.600 124.100 17.000 ;
        RECT 123.800 16.100 124.100 16.600 ;
        RECT 124.900 16.500 126.000 16.800 ;
        RECT 124.900 16.400 125.300 16.500 ;
        RECT 123.800 15.800 125.000 16.100 ;
        RECT 121.400 15.300 123.500 15.600 ;
        RECT 121.400 13.600 121.800 15.300 ;
        RECT 123.100 15.200 123.500 15.300 ;
        RECT 124.700 15.200 125.000 15.800 ;
        RECT 125.700 15.900 126.000 16.500 ;
        RECT 126.300 16.500 126.700 16.600 ;
        RECT 128.600 16.500 129.000 16.600 ;
        RECT 126.300 16.200 129.000 16.500 ;
        RECT 125.700 15.700 128.100 15.900 ;
        RECT 130.200 15.700 130.600 19.900 ;
        RECT 132.300 16.300 132.700 19.900 ;
        RECT 131.800 15.900 132.700 16.300 ;
        RECT 133.800 16.800 134.200 17.200 ;
        RECT 133.800 16.200 134.100 16.800 ;
        RECT 134.500 16.200 134.900 19.900 ;
        RECT 133.400 15.900 134.100 16.200 ;
        RECT 134.400 15.900 134.900 16.200 ;
        RECT 137.900 16.200 138.300 19.900 ;
        RECT 138.600 16.800 139.000 17.200 ;
        RECT 138.700 16.200 139.000 16.800 ;
        RECT 139.800 16.200 140.200 19.900 ;
        RECT 141.400 16.200 141.800 19.900 ;
        RECT 137.900 15.900 138.400 16.200 ;
        RECT 138.700 15.900 139.400 16.200 ;
        RECT 139.800 15.900 141.800 16.200 ;
        RECT 142.200 15.900 142.600 19.900 ;
        RECT 125.700 15.600 130.600 15.700 ;
        RECT 127.700 15.500 130.600 15.600 ;
        RECT 127.800 15.400 130.600 15.500 ;
        RECT 122.300 14.900 122.700 15.000 ;
        RECT 122.300 14.600 124.200 14.900 ;
        RECT 124.600 14.800 125.000 15.200 ;
        RECT 127.000 15.100 127.400 15.200 ;
        RECT 127.000 14.800 129.500 15.100 ;
        RECT 123.800 14.500 124.200 14.600 ;
        RECT 124.700 14.200 125.000 14.800 ;
        RECT 127.800 14.700 128.200 14.800 ;
        RECT 129.100 14.700 129.500 14.800 ;
        RECT 128.300 14.200 128.700 14.300 ;
        RECT 131.900 14.200 132.200 15.900 ;
        RECT 133.400 15.800 133.800 15.900 ;
        RECT 132.600 15.100 133.000 15.600 ;
        RECT 134.400 15.100 134.700 15.900 ;
        RECT 132.600 14.800 134.700 15.100 ;
        RECT 134.400 14.200 134.700 14.800 ;
        RECT 135.000 14.400 135.400 15.200 ;
        RECT 137.400 14.400 137.800 15.200 ;
        RECT 138.100 14.200 138.400 15.900 ;
        RECT 139.000 15.800 139.400 15.900 ;
        RECT 140.200 15.200 140.600 15.400 ;
        RECT 142.200 15.200 142.500 15.900 ;
        RECT 143.000 15.700 143.400 19.900 ;
        RECT 145.200 18.200 145.600 19.900 ;
        RECT 144.600 17.900 145.600 18.200 ;
        RECT 147.400 17.900 147.800 19.900 ;
        RECT 149.500 17.900 150.100 19.900 ;
        RECT 151.800 19.100 152.200 19.900 ;
        RECT 152.600 19.100 153.000 19.200 ;
        RECT 151.800 18.800 153.000 19.100 ;
        RECT 144.600 17.500 145.000 17.900 ;
        RECT 147.400 17.600 147.700 17.900 ;
        RECT 146.300 17.300 148.100 17.600 ;
        RECT 149.400 17.500 149.800 17.900 ;
        RECT 146.300 17.200 146.700 17.300 ;
        RECT 147.700 17.200 148.100 17.300 ;
        RECT 149.900 17.000 150.600 17.200 ;
        RECT 149.500 16.800 150.600 17.000 ;
        RECT 144.600 16.500 145.000 16.600 ;
        RECT 146.900 16.500 147.300 16.600 ;
        RECT 144.600 16.200 147.300 16.500 ;
        RECT 147.600 16.500 148.700 16.800 ;
        RECT 147.600 15.900 147.900 16.500 ;
        RECT 148.300 16.400 148.700 16.500 ;
        RECT 149.500 16.600 150.200 16.800 ;
        RECT 149.500 16.100 149.800 16.600 ;
        RECT 145.500 15.700 147.900 15.900 ;
        RECT 143.000 15.600 147.900 15.700 ;
        RECT 148.600 15.800 149.800 16.100 ;
        RECT 143.000 15.500 145.900 15.600 ;
        RECT 143.000 15.400 145.800 15.500 ;
        RECT 139.000 14.800 139.400 15.200 ;
        RECT 139.800 14.900 140.600 15.200 ;
        RECT 141.400 14.900 142.600 15.200 ;
        RECT 146.200 15.100 146.600 15.200 ;
        RECT 139.800 14.800 140.200 14.900 ;
        RECT 139.000 14.200 139.300 14.800 ;
        RECT 124.700 13.900 130.200 14.200 ;
        RECT 124.900 13.800 125.300 13.900 ;
        RECT 121.400 13.300 123.400 13.600 ;
        RECT 119.000 12.800 120.200 13.100 ;
        RECT 119.000 12.400 119.400 12.800 ;
        RECT 118.200 11.100 118.600 12.100 ;
        RECT 119.800 11.100 120.200 12.800 ;
        RECT 120.600 13.100 121.000 13.200 ;
        RECT 121.400 13.100 121.800 13.300 ;
        RECT 122.900 13.200 123.400 13.300 ;
        RECT 120.600 12.800 121.800 13.100 ;
        RECT 123.000 12.800 123.400 13.200 ;
        RECT 127.800 12.800 128.100 13.900 ;
        RECT 129.400 13.800 130.200 13.900 ;
        RECT 131.800 13.800 132.200 14.200 ;
        RECT 133.400 13.800 134.700 14.200 ;
        RECT 135.800 14.100 136.200 14.200 ;
        RECT 135.400 13.800 136.200 14.100 ;
        RECT 136.600 14.100 137.000 14.200 ;
        RECT 136.600 13.800 137.400 14.100 ;
        RECT 138.100 13.800 139.400 14.200 ;
        RECT 140.600 13.800 141.000 14.600 ;
        RECT 120.600 12.400 121.000 12.800 ;
        RECT 121.400 11.100 121.800 12.800 ;
        RECT 126.900 12.700 127.300 12.800 ;
        RECT 123.800 12.100 124.200 12.500 ;
        RECT 125.900 12.400 127.300 12.700 ;
        RECT 127.800 12.400 128.200 12.800 ;
        RECT 125.900 12.100 126.200 12.400 ;
        RECT 128.600 12.100 129.000 12.500 ;
        RECT 123.500 11.800 124.200 12.100 ;
        RECT 123.500 11.100 124.100 11.800 ;
        RECT 125.800 11.100 126.200 12.100 ;
        RECT 128.000 11.800 129.000 12.100 ;
        RECT 128.000 11.100 128.400 11.800 ;
        RECT 130.200 11.100 130.600 13.500 ;
        RECT 131.000 12.400 131.400 13.200 ;
        RECT 131.900 12.200 132.200 13.800 ;
        RECT 133.500 13.100 133.800 13.800 ;
        RECT 135.400 13.600 135.800 13.800 ;
        RECT 137.000 13.600 137.400 13.800 ;
        RECT 134.300 13.100 136.100 13.300 ;
        RECT 136.700 13.100 138.500 13.300 ;
        RECT 139.000 13.100 139.300 13.800 ;
        RECT 141.400 13.100 141.700 14.900 ;
        RECT 142.200 14.800 142.600 14.900 ;
        RECT 144.100 14.800 146.600 15.100 ;
        RECT 144.100 14.700 144.500 14.800 ;
        RECT 145.400 14.700 145.800 14.800 ;
        RECT 144.900 14.200 145.300 14.300 ;
        RECT 148.600 14.200 148.900 15.800 ;
        RECT 151.800 15.600 152.200 18.800 ;
        RECT 150.100 15.300 152.200 15.600 ;
        RECT 150.100 15.200 150.500 15.300 ;
        RECT 150.900 14.900 151.300 15.000 ;
        RECT 149.400 14.600 151.300 14.900 ;
        RECT 149.400 14.500 149.800 14.600 ;
        RECT 143.400 13.900 148.900 14.200 ;
        RECT 143.400 13.800 144.200 13.900 ;
        RECT 131.800 11.100 132.200 12.200 ;
        RECT 133.400 11.100 133.800 13.100 ;
        RECT 134.200 13.000 136.200 13.100 ;
        RECT 134.200 11.100 134.600 13.000 ;
        RECT 135.800 11.100 136.200 13.000 ;
        RECT 136.600 13.000 138.600 13.100 ;
        RECT 136.600 11.100 137.000 13.000 ;
        RECT 138.200 11.100 138.600 13.000 ;
        RECT 139.000 11.100 139.400 13.100 ;
        RECT 141.400 11.100 141.800 13.100 ;
        RECT 142.200 12.800 142.600 13.200 ;
        RECT 142.100 12.400 142.500 12.800 ;
        RECT 143.000 11.100 143.400 13.500 ;
        RECT 145.500 13.200 145.800 13.900 ;
        RECT 148.300 13.800 148.700 13.900 ;
        RECT 151.800 13.600 152.200 15.300 ;
        RECT 150.300 13.300 152.200 13.600 ;
        RECT 154.200 13.400 154.600 14.200 ;
        RECT 150.300 13.200 150.700 13.300 ;
        RECT 144.600 12.100 145.000 12.500 ;
        RECT 145.400 12.400 145.800 13.200 ;
        RECT 146.300 12.700 146.700 12.800 ;
        RECT 146.300 12.400 147.700 12.700 ;
        RECT 147.400 12.100 147.700 12.400 ;
        RECT 149.400 12.100 149.800 12.500 ;
        RECT 144.600 11.800 145.600 12.100 ;
        RECT 145.200 11.100 145.600 11.800 ;
        RECT 147.400 11.100 147.800 12.100 ;
        RECT 149.400 11.800 150.100 12.100 ;
        RECT 149.500 11.100 150.100 11.800 ;
        RECT 151.800 11.100 152.200 13.300 ;
        RECT 155.000 11.100 155.400 19.900 ;
        RECT 156.100 16.200 156.500 19.900 ;
        RECT 155.800 15.900 156.500 16.200 ;
        RECT 155.800 15.200 156.100 15.900 ;
        RECT 158.200 15.600 158.600 19.900 ;
        RECT 156.600 15.400 158.600 15.600 ;
        RECT 159.000 15.700 159.400 19.900 ;
        RECT 161.200 18.200 161.600 19.900 ;
        RECT 160.600 17.900 161.600 18.200 ;
        RECT 163.400 17.900 163.800 19.900 ;
        RECT 165.500 17.900 166.100 19.900 ;
        RECT 160.600 17.500 161.000 17.900 ;
        RECT 163.400 17.600 163.700 17.900 ;
        RECT 162.300 17.300 164.100 17.600 ;
        RECT 165.400 17.500 165.800 17.900 ;
        RECT 162.300 17.200 162.700 17.300 ;
        RECT 163.700 17.200 164.100 17.300 ;
        RECT 160.600 16.500 161.000 16.600 ;
        RECT 162.900 16.500 163.300 16.600 ;
        RECT 160.600 16.200 163.300 16.500 ;
        RECT 163.600 16.500 164.700 16.800 ;
        RECT 163.600 15.900 163.900 16.500 ;
        RECT 164.300 16.400 164.700 16.500 ;
        RECT 165.500 16.600 166.200 17.000 ;
        RECT 165.500 16.100 165.800 16.600 ;
        RECT 161.500 15.700 163.900 15.900 ;
        RECT 159.000 15.600 163.900 15.700 ;
        RECT 164.600 15.800 165.800 16.100 ;
        RECT 159.000 15.500 161.900 15.600 ;
        RECT 159.000 15.400 161.800 15.500 ;
        RECT 156.500 15.300 158.600 15.400 ;
        RECT 155.800 14.800 156.200 15.200 ;
        RECT 156.500 15.000 156.900 15.300 ;
        RECT 162.200 15.100 162.600 15.200 ;
        RECT 163.000 15.100 163.400 15.200 ;
        RECT 155.800 13.100 156.100 14.800 ;
        RECT 156.500 13.500 156.800 15.000 ;
        RECT 160.100 14.800 163.400 15.100 ;
        RECT 160.100 14.700 160.500 14.800 ;
        RECT 157.200 14.200 157.600 14.600 ;
        RECT 160.900 14.200 161.300 14.300 ;
        RECT 164.600 14.200 164.900 15.800 ;
        RECT 167.800 15.600 168.200 19.900 ;
        RECT 168.600 15.800 169.000 16.600 ;
        RECT 166.100 15.300 168.200 15.600 ;
        RECT 166.100 15.200 166.500 15.300 ;
        RECT 166.900 14.900 167.300 15.000 ;
        RECT 165.400 14.600 167.300 14.900 ;
        RECT 165.400 14.500 165.800 14.600 ;
        RECT 157.300 13.800 157.800 14.200 ;
        RECT 158.200 14.100 158.600 14.200 ;
        RECT 159.400 14.100 164.900 14.200 ;
        RECT 158.200 13.900 164.900 14.100 ;
        RECT 158.200 13.800 160.200 13.900 ;
        RECT 156.500 13.200 157.700 13.500 ;
        RECT 155.800 11.100 156.200 13.100 ;
        RECT 157.400 12.100 157.700 13.200 ;
        RECT 158.200 12.400 158.600 13.200 ;
        RECT 157.400 11.100 157.800 12.100 ;
        RECT 159.000 11.100 159.400 13.500 ;
        RECT 161.500 12.800 161.800 13.900 ;
        RECT 164.300 13.800 164.700 13.900 ;
        RECT 167.800 13.600 168.200 15.300 ;
        RECT 166.300 13.300 168.200 13.600 ;
        RECT 166.300 13.200 166.700 13.300 ;
        RECT 160.600 12.100 161.000 12.500 ;
        RECT 161.400 12.400 161.800 12.800 ;
        RECT 162.300 12.700 162.700 12.800 ;
        RECT 162.300 12.400 163.700 12.700 ;
        RECT 163.400 12.100 163.700 12.400 ;
        RECT 165.400 12.100 165.800 12.500 ;
        RECT 160.600 11.800 161.600 12.100 ;
        RECT 161.200 11.100 161.600 11.800 ;
        RECT 163.400 11.100 163.800 12.100 ;
        RECT 165.400 11.800 166.100 12.100 ;
        RECT 165.500 11.100 166.100 11.800 ;
        RECT 167.800 11.100 168.200 13.300 ;
        RECT 169.400 13.100 169.800 19.900 ;
        RECT 171.000 15.900 171.400 19.900 ;
        RECT 171.800 16.200 172.200 19.900 ;
        RECT 173.400 16.200 173.800 19.900 ;
        RECT 171.800 15.900 173.800 16.200 ;
        RECT 171.100 15.200 171.400 15.900 ;
        RECT 173.000 15.200 173.400 15.400 ;
        RECT 171.000 14.900 172.200 15.200 ;
        RECT 173.000 14.900 173.800 15.200 ;
        RECT 171.000 14.800 171.400 14.900 ;
        RECT 170.200 14.100 170.600 14.200 ;
        RECT 170.200 13.800 171.300 14.100 ;
        RECT 170.200 13.400 170.600 13.800 ;
        RECT 168.900 12.800 169.800 13.100 ;
        RECT 171.000 13.200 171.300 13.800 ;
        RECT 171.000 12.800 171.400 13.200 ;
        RECT 171.900 13.100 172.200 14.900 ;
        RECT 173.400 14.800 173.800 14.900 ;
        RECT 172.600 14.100 173.000 14.600 ;
        RECT 174.200 14.100 174.600 19.900 ;
        RECT 175.800 15.800 176.200 16.600 ;
        RECT 172.600 13.800 174.600 14.100 ;
        RECT 168.900 12.200 169.300 12.800 ;
        RECT 171.100 12.400 171.500 12.800 ;
        RECT 168.600 11.800 169.300 12.200 ;
        RECT 168.900 11.100 169.300 11.800 ;
        RECT 171.800 11.100 172.200 13.100 ;
        RECT 174.200 11.100 174.600 13.800 ;
        RECT 175.000 14.100 175.400 14.200 ;
        RECT 176.600 14.100 177.000 19.900 ;
        RECT 178.600 16.800 179.000 17.200 ;
        RECT 178.600 16.200 178.900 16.800 ;
        RECT 179.300 16.200 179.700 19.900 ;
        RECT 178.200 15.900 178.900 16.200 ;
        RECT 179.200 15.900 179.700 16.200 ;
        RECT 181.700 16.300 182.100 19.900 ;
        RECT 181.700 15.900 182.600 16.300 ;
        RECT 178.200 15.800 178.600 15.900 ;
        RECT 179.200 15.200 179.500 15.900 ;
        RECT 179.000 14.800 179.500 15.200 ;
        RECT 179.200 14.200 179.500 14.800 ;
        RECT 179.800 14.400 180.200 15.200 ;
        RECT 181.400 14.800 181.800 15.600 ;
        RECT 182.200 15.100 182.500 15.900 ;
        RECT 183.000 15.100 183.400 15.200 ;
        RECT 182.200 14.800 183.400 15.100 ;
        RECT 182.200 14.200 182.500 14.800 ;
        RECT 175.000 13.800 177.000 14.100 ;
        RECT 175.000 13.400 175.400 13.800 ;
        RECT 176.600 13.100 177.000 13.800 ;
        RECT 177.400 13.400 177.800 14.200 ;
        RECT 178.200 13.800 179.500 14.200 ;
        RECT 180.600 14.100 181.000 14.200 ;
        RECT 180.200 13.800 181.000 14.100 ;
        RECT 182.200 13.800 182.600 14.200 ;
        RECT 178.300 13.100 178.600 13.800 ;
        RECT 180.200 13.600 180.600 13.800 ;
        RECT 179.100 13.100 180.900 13.300 ;
        RECT 176.100 12.800 177.000 13.100 ;
        RECT 176.100 12.200 176.500 12.800 ;
        RECT 175.800 11.800 176.500 12.200 ;
        RECT 176.100 11.100 176.500 11.800 ;
        RECT 178.200 11.100 178.600 13.100 ;
        RECT 179.000 13.000 181.000 13.100 ;
        RECT 179.000 11.100 179.400 13.000 ;
        RECT 180.600 11.100 181.000 13.000 ;
        RECT 182.200 12.100 182.500 13.800 ;
        RECT 183.000 12.400 183.400 13.200 ;
        RECT 183.800 12.400 184.200 13.200 ;
        RECT 182.200 11.100 182.600 12.100 ;
        RECT 184.600 11.100 185.000 19.900 ;
        RECT 185.400 15.700 185.800 19.900 ;
        RECT 187.600 18.200 188.000 19.900 ;
        RECT 187.000 17.900 188.000 18.200 ;
        RECT 189.800 17.900 190.200 19.900 ;
        RECT 191.900 17.900 192.500 19.900 ;
        RECT 187.000 17.500 187.400 17.900 ;
        RECT 189.800 17.600 190.100 17.900 ;
        RECT 188.700 17.300 190.500 17.600 ;
        RECT 191.800 17.500 192.200 17.900 ;
        RECT 188.700 17.200 189.100 17.300 ;
        RECT 190.100 17.200 190.500 17.300 ;
        RECT 187.000 16.500 187.400 16.600 ;
        RECT 189.300 16.500 189.700 16.600 ;
        RECT 187.000 16.200 189.700 16.500 ;
        RECT 190.000 16.500 191.100 16.800 ;
        RECT 190.000 15.900 190.300 16.500 ;
        RECT 190.700 16.400 191.100 16.500 ;
        RECT 191.900 16.600 192.600 17.000 ;
        RECT 191.900 16.100 192.200 16.600 ;
        RECT 187.900 15.700 190.300 15.900 ;
        RECT 185.400 15.600 190.300 15.700 ;
        RECT 191.000 15.800 192.200 16.100 ;
        RECT 185.400 15.500 188.300 15.600 ;
        RECT 185.400 15.400 188.200 15.500 ;
        RECT 188.600 15.100 189.000 15.200 ;
        RECT 186.500 14.800 189.000 15.100 ;
        RECT 186.500 14.700 186.900 14.800 ;
        RECT 187.800 14.700 188.200 14.800 ;
        RECT 187.300 14.200 187.700 14.300 ;
        RECT 191.000 14.200 191.300 15.800 ;
        RECT 194.200 15.600 194.600 19.900 ;
        RECT 192.500 15.300 194.600 15.600 ;
        RECT 192.500 15.200 192.900 15.300 ;
        RECT 193.300 14.900 193.700 15.000 ;
        RECT 191.800 14.600 193.700 14.900 ;
        RECT 191.800 14.500 192.200 14.600 ;
        RECT 185.800 13.900 191.300 14.200 ;
        RECT 185.800 13.800 186.600 13.900 ;
        RECT 185.400 11.100 185.800 13.500 ;
        RECT 187.900 12.800 188.200 13.900 ;
        RECT 190.700 13.800 191.100 13.900 ;
        RECT 194.200 13.600 194.600 15.300 ;
        RECT 192.700 13.300 194.600 13.600 ;
        RECT 192.700 13.200 193.100 13.300 ;
        RECT 187.000 12.100 187.400 12.500 ;
        RECT 187.800 12.400 188.200 12.800 ;
        RECT 188.700 12.700 189.100 12.800 ;
        RECT 188.700 12.400 190.100 12.700 ;
        RECT 189.800 12.100 190.100 12.400 ;
        RECT 191.800 12.100 192.200 12.500 ;
        RECT 187.000 11.800 188.000 12.100 ;
        RECT 187.600 11.100 188.000 11.800 ;
        RECT 189.800 11.100 190.200 12.100 ;
        RECT 191.800 11.800 192.500 12.100 ;
        RECT 191.900 11.100 192.500 11.800 ;
        RECT 194.200 11.100 194.600 13.300 ;
        RECT 0.600 7.800 1.000 8.600 ;
        RECT 1.400 7.100 1.800 9.900 ;
        RECT 2.200 8.000 2.600 9.900 ;
        RECT 3.800 8.000 4.200 9.900 ;
        RECT 2.200 7.900 4.200 8.000 ;
        RECT 4.600 7.900 5.000 9.900 ;
        RECT 6.200 8.900 6.600 9.900 ;
        RECT 10.200 8.900 10.600 9.900 ;
        RECT 11.800 9.200 12.200 9.900 ;
        RECT 2.300 7.700 4.100 7.900 ;
        RECT 2.600 7.200 3.000 7.400 ;
        RECT 4.600 7.200 4.900 7.900 ;
        RECT 6.200 7.200 6.500 8.900 ;
        RECT 10.000 8.800 10.600 8.900 ;
        RECT 11.700 8.800 12.200 9.200 ;
        RECT 15.000 8.900 15.400 9.900 ;
        RECT 7.000 7.800 7.400 8.600 ;
        RECT 10.000 8.500 12.000 8.800 ;
        RECT 2.200 7.100 3.000 7.200 ;
        RECT 1.400 6.900 3.000 7.100 ;
        RECT 1.400 6.800 2.600 6.900 ;
        RECT 3.700 6.800 5.000 7.200 ;
        RECT 6.200 7.100 6.600 7.200 ;
        RECT 8.600 7.100 9.000 7.200 ;
        RECT 6.200 6.800 9.000 7.100 ;
        RECT 1.400 1.100 1.800 6.800 ;
        RECT 3.000 5.800 3.400 6.600 ;
        RECT 3.700 6.100 4.000 6.800 ;
        RECT 5.400 6.100 5.800 6.200 ;
        RECT 3.700 5.800 5.800 6.100 ;
        RECT 3.700 5.100 4.000 5.800 ;
        RECT 5.400 5.400 5.800 5.800 ;
        RECT 4.600 5.100 5.000 5.200 ;
        RECT 6.200 5.100 6.500 6.800 ;
        RECT 10.000 5.200 10.300 8.500 ;
        RECT 12.100 7.800 13.000 8.200 ;
        RECT 15.000 7.200 15.300 8.900 ;
        RECT 15.800 7.800 16.200 8.600 ;
        RECT 16.900 8.200 17.300 9.900 ;
        RECT 16.900 7.900 17.800 8.200 ;
        RECT 19.000 7.900 19.400 9.900 ;
        RECT 19.800 8.000 20.200 9.900 ;
        RECT 21.400 8.000 21.800 9.900 ;
        RECT 19.800 7.900 21.800 8.000 ;
        RECT 23.000 8.100 23.400 9.900 ;
        RECT 24.600 8.900 25.000 9.900 ;
        RECT 28.600 8.900 29.000 9.900 ;
        RECT 30.200 9.200 30.600 9.900 ;
        RECT 23.800 8.100 24.200 8.600 ;
        RECT 24.700 8.100 25.000 8.900 ;
        RECT 28.400 8.800 29.000 8.900 ;
        RECT 30.100 8.800 30.600 9.200 ;
        RECT 32.900 9.200 33.300 9.900 ;
        RECT 32.900 8.800 33.800 9.200 ;
        RECT 28.400 8.500 30.400 8.800 ;
        RECT 27.000 8.100 27.400 8.200 ;
        RECT 11.400 6.800 12.200 7.200 ;
        RECT 15.000 7.100 15.400 7.200 ;
        RECT 12.600 6.800 15.400 7.100 ;
        RECT 10.600 6.100 11.400 6.200 ;
        RECT 12.600 6.100 12.900 6.800 ;
        RECT 10.600 5.800 12.900 6.100 ;
        RECT 14.200 5.400 14.600 6.200 ;
        RECT 3.500 4.800 4.000 5.100 ;
        RECT 4.300 4.800 5.000 5.100 ;
        RECT 3.500 1.100 3.900 4.800 ;
        RECT 4.300 4.200 4.600 4.800 ;
        RECT 4.200 3.800 4.600 4.200 ;
        RECT 5.700 4.700 6.600 5.100 ;
        RECT 8.600 4.900 10.300 5.200 ;
        RECT 15.000 5.100 15.300 6.800 ;
        RECT 15.800 6.100 16.200 6.200 ;
        RECT 17.400 6.100 17.800 7.900 ;
        RECT 18.200 6.800 18.600 7.600 ;
        RECT 19.100 7.200 19.400 7.900 ;
        RECT 19.900 7.700 21.700 7.900 ;
        RECT 23.000 7.800 24.200 8.100 ;
        RECT 24.600 7.800 27.400 8.100 ;
        RECT 21.000 7.200 21.400 7.400 ;
        RECT 19.000 6.800 20.300 7.200 ;
        RECT 21.000 6.900 21.800 7.200 ;
        RECT 21.400 6.800 21.800 6.900 ;
        RECT 22.200 6.800 22.600 7.600 ;
        RECT 15.800 5.800 17.800 6.100 ;
        RECT 8.600 4.800 9.000 4.900 ;
        RECT 5.700 1.100 6.100 4.700 ;
        RECT 8.700 4.500 9.000 4.800 ;
        RECT 14.500 4.700 15.400 5.100 ;
        RECT 9.500 4.500 11.300 4.600 ;
        RECT 7.800 1.500 8.200 4.500 ;
        RECT 8.600 1.700 9.000 4.500 ;
        RECT 9.400 4.300 11.300 4.500 ;
        RECT 7.900 1.400 8.200 1.500 ;
        RECT 9.400 1.500 9.800 4.300 ;
        RECT 11.000 4.100 11.300 4.300 ;
        RECT 11.900 4.400 13.700 4.700 ;
        RECT 11.900 4.100 12.200 4.400 ;
        RECT 9.400 1.400 9.700 1.500 ;
        RECT 7.900 1.100 9.700 1.400 ;
        RECT 10.200 1.400 10.600 4.000 ;
        RECT 11.000 1.700 11.400 4.100 ;
        RECT 11.800 1.400 12.200 4.100 ;
        RECT 10.200 1.100 12.200 1.400 ;
        RECT 13.400 4.100 13.700 4.400 ;
        RECT 13.400 1.100 13.800 4.100 ;
        RECT 14.500 1.100 14.900 4.700 ;
        RECT 16.600 4.400 17.000 5.200 ;
        RECT 17.400 1.100 17.800 5.800 ;
        RECT 19.000 5.100 19.400 5.200 ;
        RECT 20.000 5.100 20.300 6.800 ;
        RECT 20.600 5.800 21.000 6.600 ;
        RECT 19.000 4.800 19.700 5.100 ;
        RECT 20.000 4.800 20.500 5.100 ;
        RECT 19.400 4.200 19.700 4.800 ;
        RECT 19.400 3.800 19.800 4.200 ;
        RECT 20.100 1.100 20.500 4.800 ;
        RECT 23.000 1.100 23.400 7.800 ;
        RECT 23.800 7.200 24.100 7.800 ;
        RECT 24.700 7.200 25.000 7.800 ;
        RECT 23.800 6.800 24.200 7.200 ;
        RECT 24.600 6.800 25.000 7.200 ;
        RECT 24.700 5.100 25.000 6.800 ;
        RECT 25.400 5.400 25.800 6.200 ;
        RECT 28.400 5.200 28.700 8.500 ;
        RECT 32.900 8.200 33.300 8.800 ;
        RECT 30.200 7.800 31.400 8.200 ;
        RECT 32.900 7.900 33.800 8.200 ;
        RECT 29.800 7.100 30.600 7.200 ;
        RECT 31.000 7.100 31.400 7.200 ;
        RECT 29.800 6.800 31.400 7.100 ;
        RECT 29.000 5.800 29.800 6.200 ;
        RECT 24.600 4.700 25.500 5.100 ;
        RECT 27.000 4.900 28.700 5.200 ;
        RECT 27.000 4.800 27.400 4.900 ;
        RECT 25.100 1.100 25.500 4.700 ;
        RECT 27.100 4.500 27.400 4.800 ;
        RECT 27.900 4.500 29.700 4.600 ;
        RECT 26.200 1.500 26.600 4.500 ;
        RECT 27.000 1.700 27.400 4.500 ;
        RECT 27.800 4.300 29.700 4.500 ;
        RECT 26.300 1.400 26.600 1.500 ;
        RECT 27.800 1.500 28.200 4.300 ;
        RECT 29.400 4.100 29.700 4.300 ;
        RECT 30.300 4.400 32.100 4.700 ;
        RECT 32.600 4.400 33.000 5.200 ;
        RECT 30.300 4.100 30.600 4.400 ;
        RECT 27.800 1.400 28.100 1.500 ;
        RECT 26.300 1.100 28.100 1.400 ;
        RECT 28.600 1.400 29.000 4.000 ;
        RECT 29.400 1.700 29.800 4.100 ;
        RECT 30.200 1.400 30.600 4.100 ;
        RECT 28.600 1.100 30.600 1.400 ;
        RECT 31.800 4.100 32.100 4.400 ;
        RECT 31.800 1.100 32.200 4.100 ;
        RECT 33.400 1.100 33.800 7.900 ;
        RECT 35.000 7.700 35.400 9.900 ;
        RECT 37.100 9.200 37.700 9.900 ;
        RECT 37.100 8.900 37.800 9.200 ;
        RECT 39.400 8.900 39.800 9.900 ;
        RECT 41.600 9.200 42.000 9.900 ;
        RECT 41.600 8.900 42.600 9.200 ;
        RECT 37.400 8.500 37.800 8.900 ;
        RECT 39.500 8.600 39.800 8.900 ;
        RECT 39.500 8.300 40.900 8.600 ;
        RECT 40.500 8.200 40.900 8.300 ;
        RECT 41.400 7.800 41.800 8.600 ;
        RECT 42.200 8.500 42.600 8.900 ;
        RECT 36.500 7.700 36.900 7.800 ;
        RECT 34.200 7.100 34.600 7.600 ;
        RECT 35.000 7.400 36.900 7.700 ;
        RECT 35.000 7.100 35.400 7.400 ;
        RECT 38.500 7.100 38.900 7.200 ;
        RECT 41.400 7.100 41.700 7.800 ;
        RECT 43.800 7.500 44.200 9.900 ;
        RECT 46.200 8.000 46.600 9.900 ;
        RECT 47.800 8.000 48.200 9.900 ;
        RECT 46.200 7.900 48.200 8.000 ;
        RECT 48.600 7.900 49.000 9.900 ;
        RECT 50.200 8.800 50.600 9.900 ;
        RECT 46.300 7.700 48.100 7.900 ;
        RECT 46.600 7.200 47.000 7.400 ;
        RECT 48.600 7.200 48.900 7.900 ;
        RECT 49.400 7.800 49.800 8.600 ;
        RECT 50.300 7.200 50.600 8.800 ;
        RECT 51.800 7.800 52.200 8.600 ;
        RECT 43.000 7.100 43.800 7.200 ;
        RECT 34.200 6.800 35.400 7.100 ;
        RECT 35.000 5.700 35.400 6.800 ;
        RECT 38.300 6.800 43.800 7.100 ;
        RECT 46.200 6.900 47.000 7.200 ;
        RECT 46.200 6.800 46.600 6.900 ;
        RECT 47.700 6.800 49.000 7.200 ;
        RECT 50.200 6.800 50.600 7.200 ;
        RECT 37.400 6.400 37.800 6.500 ;
        RECT 35.900 6.100 37.800 6.400 ;
        RECT 35.900 6.000 36.300 6.100 ;
        RECT 36.700 5.700 37.100 5.800 ;
        RECT 35.000 5.400 37.100 5.700 ;
        RECT 35.000 1.100 35.400 5.400 ;
        RECT 38.300 5.200 38.600 6.800 ;
        RECT 41.900 6.700 42.300 6.800 ;
        RECT 41.400 6.200 41.800 6.300 ;
        RECT 42.700 6.200 43.100 6.300 ;
        RECT 40.600 5.900 43.100 6.200 ;
        RECT 45.400 6.100 45.800 6.200 ;
        RECT 47.000 6.100 47.400 6.600 ;
        RECT 40.600 5.800 41.000 5.900 ;
        RECT 45.400 5.800 47.400 6.100 ;
        RECT 47.700 6.100 48.000 6.800 ;
        RECT 49.400 6.100 49.800 6.200 ;
        RECT 47.700 5.800 49.800 6.100 ;
        RECT 41.400 5.500 44.200 5.600 ;
        RECT 41.300 5.400 44.200 5.500 ;
        RECT 37.400 4.900 38.600 5.200 ;
        RECT 39.300 5.300 44.200 5.400 ;
        RECT 39.300 5.100 41.700 5.300 ;
        RECT 37.400 4.400 37.700 4.900 ;
        RECT 37.000 4.000 37.700 4.400 ;
        RECT 38.500 4.500 38.900 4.600 ;
        RECT 39.300 4.500 39.600 5.100 ;
        RECT 38.500 4.200 39.600 4.500 ;
        RECT 39.900 4.500 42.600 4.800 ;
        RECT 39.900 4.400 40.300 4.500 ;
        RECT 42.200 4.400 42.600 4.500 ;
        RECT 39.100 3.700 39.500 3.800 ;
        RECT 40.500 3.700 40.900 3.800 ;
        RECT 37.400 3.100 37.800 3.500 ;
        RECT 39.100 3.400 40.900 3.700 ;
        RECT 39.500 3.100 39.800 3.400 ;
        RECT 42.200 3.100 42.600 3.500 ;
        RECT 37.100 1.100 37.700 3.100 ;
        RECT 39.400 1.100 39.800 3.100 ;
        RECT 41.600 2.800 42.600 3.100 ;
        RECT 41.600 1.100 42.000 2.800 ;
        RECT 43.800 1.100 44.200 5.300 ;
        RECT 47.700 5.100 48.000 5.800 ;
        RECT 48.600 5.100 49.000 5.200 ;
        RECT 50.300 5.100 50.600 6.800 ;
        RECT 52.600 7.100 53.000 9.900 ;
        RECT 53.400 8.000 53.800 9.900 ;
        RECT 55.000 8.000 55.400 9.900 ;
        RECT 53.400 7.900 55.400 8.000 ;
        RECT 55.800 7.900 56.200 9.900 ;
        RECT 53.500 7.700 55.300 7.900 ;
        RECT 53.800 7.200 54.200 7.400 ;
        RECT 55.800 7.200 56.100 7.900 ;
        RECT 56.600 7.600 57.000 9.900 ;
        RECT 60.600 7.800 61.000 9.900 ;
        RECT 63.500 9.200 63.900 9.900 ;
        RECT 63.500 8.800 64.200 9.200 ;
        RECT 61.300 8.200 61.700 8.600 ;
        RECT 63.500 8.200 63.900 8.800 ;
        RECT 61.400 7.800 61.800 8.200 ;
        RECT 63.000 7.900 63.900 8.200 ;
        RECT 56.600 7.300 57.700 7.600 ;
        RECT 53.400 7.100 54.200 7.200 ;
        RECT 52.600 6.900 54.200 7.100 ;
        RECT 52.600 6.800 53.800 6.900 ;
        RECT 54.900 6.800 56.200 7.200 ;
        RECT 51.000 5.400 51.400 6.200 ;
        RECT 47.500 4.800 48.000 5.100 ;
        RECT 48.300 4.800 49.000 5.100 ;
        RECT 47.500 1.100 47.900 4.800 ;
        RECT 48.300 4.200 48.600 4.800 ;
        RECT 50.200 4.700 51.100 5.100 ;
        RECT 48.200 3.800 48.600 4.200 ;
        RECT 50.700 1.100 51.100 4.700 ;
        RECT 52.600 1.100 53.000 6.800 ;
        RECT 53.400 6.100 53.800 6.200 ;
        RECT 54.200 6.100 54.600 6.600 ;
        RECT 53.400 5.800 54.600 6.100 ;
        RECT 54.900 5.200 55.200 6.800 ;
        RECT 57.400 5.800 57.700 7.300 ;
        RECT 59.800 6.400 60.200 7.200 ;
        RECT 59.000 6.100 59.400 6.200 ;
        RECT 60.600 6.100 60.900 7.800 ;
        RECT 62.200 6.800 62.600 7.600 ;
        RECT 61.400 6.100 61.800 6.200 ;
        RECT 59.000 5.800 59.800 6.100 ;
        RECT 60.600 5.800 61.800 6.100 ;
        RECT 57.400 5.400 58.000 5.800 ;
        RECT 59.400 5.600 59.800 5.800 ;
        RECT 54.200 4.800 55.200 5.200 ;
        RECT 55.800 5.100 56.200 5.200 ;
        RECT 57.400 5.100 57.700 5.400 ;
        RECT 61.400 5.100 61.700 5.800 ;
        RECT 55.500 4.800 56.200 5.100 ;
        RECT 56.600 4.800 57.700 5.100 ;
        RECT 59.000 4.800 61.000 5.100 ;
        RECT 54.700 1.100 55.100 4.800 ;
        RECT 55.500 4.200 55.800 4.800 ;
        RECT 55.400 3.800 55.800 4.200 ;
        RECT 56.600 1.100 57.000 4.800 ;
        RECT 59.000 1.100 59.400 4.800 ;
        RECT 60.600 1.100 61.000 4.800 ;
        RECT 61.400 1.100 61.800 5.100 ;
        RECT 63.000 1.100 63.400 7.900 ;
        RECT 64.600 7.500 65.000 9.900 ;
        RECT 66.800 9.200 67.200 9.900 ;
        RECT 66.200 8.900 67.200 9.200 ;
        RECT 69.000 8.900 69.400 9.900 ;
        RECT 71.100 9.200 71.700 9.900 ;
        RECT 71.000 8.900 71.700 9.200 ;
        RECT 66.200 8.500 66.600 8.900 ;
        RECT 69.000 8.600 69.300 8.900 ;
        RECT 67.000 7.800 67.400 8.600 ;
        RECT 67.900 8.300 69.300 8.600 ;
        RECT 71.000 8.500 71.400 8.900 ;
        RECT 67.900 8.200 68.300 8.300 ;
        RECT 73.400 8.100 73.800 9.900 ;
        RECT 74.200 8.100 74.600 8.600 ;
        RECT 73.400 7.800 74.600 8.100 ;
        RECT 65.000 7.100 65.800 7.200 ;
        RECT 67.100 7.100 67.400 7.800 ;
        RECT 71.900 7.700 72.300 7.800 ;
        RECT 73.400 7.700 73.800 7.800 ;
        RECT 71.900 7.400 73.800 7.700 ;
        RECT 69.900 7.100 70.300 7.200 ;
        RECT 65.000 6.800 70.500 7.100 ;
        RECT 66.500 6.700 66.900 6.800 ;
        RECT 65.700 6.200 66.100 6.300 ;
        RECT 65.700 6.100 68.200 6.200 ;
        RECT 69.400 6.100 69.800 6.200 ;
        RECT 65.700 5.900 69.800 6.100 ;
        RECT 67.800 5.800 69.800 5.900 ;
        RECT 64.600 5.500 67.400 5.600 ;
        RECT 64.600 5.400 67.500 5.500 ;
        RECT 64.600 5.300 69.500 5.400 ;
        RECT 63.800 4.400 64.200 5.200 ;
        RECT 64.600 1.100 65.000 5.300 ;
        RECT 67.100 5.100 69.500 5.300 ;
        RECT 66.200 4.500 68.900 4.800 ;
        RECT 66.200 4.400 66.600 4.500 ;
        RECT 68.500 4.400 68.900 4.500 ;
        RECT 69.200 4.500 69.500 5.100 ;
        RECT 70.200 5.200 70.500 6.800 ;
        RECT 71.000 6.400 71.400 6.500 ;
        RECT 71.000 6.100 72.900 6.400 ;
        RECT 72.500 6.000 72.900 6.100 ;
        RECT 71.700 5.700 72.100 5.800 ;
        RECT 73.400 5.700 73.800 7.400 ;
        RECT 71.700 5.400 73.800 5.700 ;
        RECT 70.200 4.900 71.400 5.200 ;
        RECT 69.900 4.500 70.300 4.600 ;
        RECT 69.200 4.200 70.300 4.500 ;
        RECT 71.100 4.400 71.400 4.900 ;
        RECT 71.100 4.000 71.800 4.400 ;
        RECT 67.900 3.700 68.300 3.800 ;
        RECT 69.300 3.700 69.700 3.800 ;
        RECT 66.200 3.100 66.600 3.500 ;
        RECT 67.900 3.400 69.700 3.700 ;
        RECT 69.000 3.100 69.300 3.400 ;
        RECT 71.000 3.100 71.400 3.500 ;
        RECT 66.200 2.800 67.200 3.100 ;
        RECT 66.800 1.100 67.200 2.800 ;
        RECT 69.000 1.100 69.400 3.100 ;
        RECT 71.100 1.100 71.700 3.100 ;
        RECT 73.400 1.100 73.800 5.400 ;
        RECT 75.000 6.100 75.400 9.900 ;
        RECT 77.400 7.900 77.800 9.900 ;
        RECT 79.800 8.900 80.200 9.900 ;
        RECT 78.100 8.200 78.500 8.600 ;
        RECT 76.600 6.400 77.000 7.200 ;
        RECT 75.800 6.100 76.200 6.200 ;
        RECT 77.400 6.100 77.700 7.900 ;
        RECT 78.200 7.800 78.600 8.200 ;
        RECT 79.000 7.800 79.400 8.600 ;
        RECT 79.900 7.800 80.200 8.900 ;
        RECT 81.400 7.900 81.800 9.900 ;
        RECT 79.900 7.500 81.100 7.800 ;
        RECT 79.800 6.800 80.300 7.200 ;
        RECT 80.000 6.400 80.400 6.800 ;
        RECT 78.200 6.100 78.600 6.200 ;
        RECT 75.000 5.800 76.600 6.100 ;
        RECT 77.400 5.800 78.600 6.100 ;
        RECT 80.800 6.000 81.100 7.500 ;
        RECT 81.500 6.200 81.800 7.900 ;
        RECT 82.200 7.800 82.600 8.600 ;
        RECT 75.000 1.100 75.400 5.800 ;
        RECT 76.200 5.600 76.600 5.800 ;
        RECT 78.200 5.100 78.500 5.800 ;
        RECT 80.700 5.700 81.100 6.000 ;
        RECT 81.400 5.800 81.800 6.200 ;
        RECT 79.000 5.600 81.100 5.700 ;
        RECT 79.000 5.400 81.000 5.600 ;
        RECT 75.800 4.800 77.800 5.100 ;
        RECT 75.800 1.100 76.200 4.800 ;
        RECT 77.400 1.100 77.800 4.800 ;
        RECT 78.200 1.100 78.600 5.100 ;
        RECT 79.000 1.100 79.400 5.400 ;
        RECT 81.500 5.100 81.800 5.800 ;
        RECT 81.100 4.800 81.800 5.100 ;
        RECT 83.000 5.100 83.400 9.900 ;
        RECT 85.600 7.100 86.000 9.900 ;
        RECT 87.300 9.200 87.700 9.900 ;
        RECT 87.000 8.800 87.700 9.200 ;
        RECT 87.300 8.200 87.700 8.800 ;
        RECT 87.300 7.900 88.200 8.200 ;
        RECT 85.600 6.900 86.500 7.100 ;
        RECT 85.700 6.800 86.500 6.900 ;
        RECT 84.600 5.800 85.800 6.200 ;
        RECT 83.800 5.100 84.200 5.600 ;
        RECT 83.000 4.800 84.200 5.100 ;
        RECT 86.200 5.200 86.500 6.800 ;
        RECT 86.200 4.800 86.600 5.200 ;
        RECT 81.100 1.100 81.500 4.800 ;
        RECT 83.000 1.100 83.400 4.800 ;
        RECT 85.400 3.800 85.800 4.600 ;
        RECT 86.200 3.500 86.500 4.800 ;
        RECT 87.000 4.400 87.400 5.200 ;
        RECT 84.700 3.200 86.500 3.500 ;
        RECT 84.600 1.100 85.000 3.200 ;
        RECT 86.200 3.100 86.500 3.200 ;
        RECT 86.200 1.100 86.600 3.100 ;
        RECT 87.800 1.100 88.200 7.900 ;
        RECT 88.600 6.800 89.000 7.600 ;
        RECT 89.400 7.500 89.800 9.900 ;
        RECT 91.600 9.200 92.000 9.900 ;
        RECT 91.000 8.900 92.000 9.200 ;
        RECT 93.800 8.900 94.200 9.900 ;
        RECT 95.900 9.200 96.500 9.900 ;
        RECT 95.800 8.900 96.500 9.200 ;
        RECT 91.000 8.500 91.400 8.900 ;
        RECT 93.800 8.600 94.100 8.900 ;
        RECT 91.800 7.800 92.200 8.600 ;
        RECT 92.700 8.300 94.100 8.600 ;
        RECT 95.800 8.500 96.200 8.900 ;
        RECT 92.700 8.200 93.100 8.300 ;
        RECT 89.800 7.100 90.600 7.200 ;
        RECT 91.900 7.100 92.200 7.800 ;
        RECT 96.700 7.700 97.100 7.800 ;
        RECT 98.200 7.700 98.600 9.900 ;
        RECT 101.400 8.900 101.800 9.900 ;
        RECT 103.300 9.200 103.700 9.900 ;
        RECT 105.700 9.200 106.100 9.900 ;
        RECT 100.600 7.800 101.000 8.600 ;
        RECT 96.700 7.400 98.600 7.700 ;
        RECT 94.700 7.100 95.100 7.200 ;
        RECT 89.800 6.800 95.300 7.100 ;
        RECT 91.300 6.700 91.700 6.800 ;
        RECT 90.500 6.200 90.900 6.300 ;
        RECT 90.500 5.900 93.000 6.200 ;
        RECT 92.600 5.800 93.000 5.900 ;
        RECT 89.400 5.500 92.200 5.600 ;
        RECT 89.400 5.400 92.300 5.500 ;
        RECT 89.400 5.300 94.300 5.400 ;
        RECT 89.400 1.100 89.800 5.300 ;
        RECT 91.900 5.100 94.300 5.300 ;
        RECT 91.000 4.500 93.700 4.800 ;
        RECT 91.000 4.400 91.400 4.500 ;
        RECT 93.300 4.400 93.700 4.500 ;
        RECT 94.000 4.500 94.300 5.100 ;
        RECT 95.000 5.200 95.300 6.800 ;
        RECT 95.800 6.400 96.200 6.500 ;
        RECT 95.800 6.100 97.700 6.400 ;
        RECT 97.300 6.000 97.700 6.100 ;
        RECT 96.500 5.700 96.900 5.800 ;
        RECT 98.200 5.700 98.600 7.400 ;
        RECT 101.500 7.200 101.800 8.900 ;
        RECT 103.000 8.800 103.700 9.200 ;
        RECT 105.400 8.800 106.100 9.200 ;
        RECT 103.300 8.200 103.700 8.800 ;
        RECT 105.700 8.400 106.100 8.800 ;
        RECT 103.300 7.900 104.200 8.200 ;
        RECT 101.400 6.800 101.800 7.200 ;
        RECT 96.500 5.400 98.600 5.700 ;
        RECT 95.000 4.900 96.200 5.200 ;
        RECT 94.700 4.500 95.100 4.600 ;
        RECT 94.000 4.200 95.100 4.500 ;
        RECT 95.900 4.400 96.200 4.900 ;
        RECT 95.900 4.000 96.600 4.400 ;
        RECT 92.700 3.700 93.100 3.800 ;
        RECT 94.100 3.700 94.500 3.800 ;
        RECT 91.000 3.100 91.400 3.500 ;
        RECT 92.700 3.400 94.500 3.700 ;
        RECT 93.800 3.100 94.100 3.400 ;
        RECT 95.800 3.100 96.200 3.500 ;
        RECT 91.000 2.800 92.000 3.100 ;
        RECT 91.600 1.100 92.000 2.800 ;
        RECT 93.800 1.100 94.200 3.100 ;
        RECT 95.900 1.100 96.500 3.100 ;
        RECT 98.200 1.100 98.600 5.400 ;
        RECT 101.500 5.100 101.800 6.800 ;
        RECT 102.200 5.400 102.600 6.200 ;
        RECT 101.400 4.700 102.300 5.100 ;
        RECT 101.900 1.100 102.300 4.700 ;
        RECT 103.000 4.400 103.400 5.200 ;
        RECT 103.800 1.100 104.200 7.900 ;
        RECT 105.400 7.900 106.100 8.400 ;
        RECT 107.800 7.900 108.200 9.900 ;
        RECT 104.600 6.800 105.000 7.600 ;
        RECT 105.400 6.200 105.700 7.900 ;
        RECT 107.800 7.800 108.100 7.900 ;
        RECT 107.200 7.600 108.100 7.800 ;
        RECT 106.000 7.500 108.100 7.600 ;
        RECT 108.600 7.700 109.000 9.900 ;
        RECT 110.700 9.200 111.300 9.900 ;
        RECT 110.700 8.900 111.400 9.200 ;
        RECT 113.000 8.900 113.400 9.900 ;
        RECT 115.200 9.200 115.600 9.900 ;
        RECT 115.200 8.900 116.200 9.200 ;
        RECT 111.000 8.500 111.400 8.900 ;
        RECT 113.100 8.600 113.400 8.900 ;
        RECT 113.100 8.300 114.500 8.600 ;
        RECT 114.100 8.200 114.500 8.300 ;
        RECT 115.000 8.200 115.400 8.600 ;
        RECT 115.800 8.500 116.200 8.900 ;
        RECT 110.100 7.700 110.500 7.800 ;
        RECT 106.000 7.300 107.500 7.500 ;
        RECT 108.600 7.400 110.500 7.700 ;
        RECT 106.000 7.200 106.400 7.300 ;
        RECT 105.400 5.800 105.800 6.200 ;
        RECT 105.400 5.100 105.700 5.800 ;
        RECT 106.100 5.500 106.400 7.200 ;
        RECT 107.800 7.100 108.200 7.200 ;
        RECT 108.600 7.100 109.000 7.400 ;
        RECT 112.100 7.100 112.500 7.200 ;
        RECT 113.400 7.100 113.800 7.200 ;
        RECT 115.000 7.100 115.300 8.200 ;
        RECT 117.400 7.500 117.800 9.900 ;
        RECT 118.500 9.200 118.900 9.900 ;
        RECT 118.200 8.800 118.900 9.200 ;
        RECT 118.500 8.200 118.900 8.800 ;
        RECT 121.400 8.900 121.800 9.900 ;
        RECT 121.400 8.200 121.700 8.900 ;
        RECT 118.500 7.900 119.400 8.200 ;
        RECT 116.600 7.100 117.400 7.200 ;
        RECT 106.800 6.900 107.200 7.000 ;
        RECT 106.800 6.600 107.300 6.900 ;
        RECT 107.000 6.200 107.300 6.600 ;
        RECT 107.800 6.800 109.000 7.100 ;
        RECT 107.800 6.400 108.200 6.800 ;
        RECT 107.000 5.800 107.400 6.200 ;
        RECT 108.600 5.700 109.000 6.800 ;
        RECT 111.900 6.800 117.400 7.100 ;
        RECT 111.000 6.400 111.400 6.500 ;
        RECT 109.500 6.100 111.400 6.400 ;
        RECT 109.500 6.000 109.900 6.100 ;
        RECT 110.300 5.700 110.700 5.800 ;
        RECT 106.100 5.200 107.300 5.500 ;
        RECT 105.400 1.100 105.800 5.100 ;
        RECT 107.000 3.100 107.300 5.200 ;
        RECT 108.600 5.400 110.700 5.700 ;
        RECT 107.000 1.100 107.400 3.100 ;
        RECT 108.600 1.100 109.000 5.400 ;
        RECT 111.900 5.200 112.200 6.800 ;
        RECT 115.500 6.700 115.900 6.800 ;
        RECT 115.000 6.200 115.400 6.300 ;
        RECT 116.300 6.200 116.700 6.300 ;
        RECT 114.200 5.900 116.700 6.200 ;
        RECT 114.200 5.800 114.600 5.900 ;
        RECT 118.200 5.800 118.600 6.200 ;
        RECT 115.000 5.500 117.800 5.600 ;
        RECT 114.900 5.400 117.800 5.500 ;
        RECT 111.000 4.900 112.200 5.200 ;
        RECT 112.900 5.300 117.800 5.400 ;
        RECT 112.900 5.100 115.300 5.300 ;
        RECT 111.000 4.400 111.300 4.900 ;
        RECT 110.600 4.000 111.300 4.400 ;
        RECT 112.100 4.500 112.500 4.600 ;
        RECT 112.900 4.500 113.200 5.100 ;
        RECT 112.100 4.200 113.200 4.500 ;
        RECT 113.500 4.500 116.200 4.800 ;
        RECT 113.500 4.400 113.900 4.500 ;
        RECT 115.800 4.400 116.200 4.500 ;
        RECT 112.700 3.700 113.100 3.800 ;
        RECT 114.100 3.700 114.500 3.800 ;
        RECT 111.000 3.100 111.400 3.500 ;
        RECT 112.700 3.400 114.500 3.700 ;
        RECT 113.100 3.100 113.400 3.400 ;
        RECT 115.800 3.100 116.200 3.500 ;
        RECT 110.700 1.100 111.300 3.100 ;
        RECT 113.000 1.100 113.400 3.100 ;
        RECT 115.200 2.800 116.200 3.100 ;
        RECT 115.200 1.100 115.600 2.800 ;
        RECT 117.400 1.100 117.800 5.300 ;
        RECT 118.200 5.200 118.500 5.800 ;
        RECT 118.200 4.400 118.600 5.200 ;
        RECT 119.000 1.100 119.400 7.900 ;
        RECT 121.400 7.800 121.800 8.200 ;
        RECT 122.200 7.800 122.600 8.600 ;
        RECT 123.000 8.000 123.400 9.900 ;
        RECT 124.600 8.000 125.000 9.900 ;
        RECT 123.000 7.900 125.000 8.000 ;
        RECT 125.400 7.900 125.800 9.900 ;
        RECT 127.500 8.200 127.900 9.900 ;
        RECT 127.000 7.900 127.900 8.200 ;
        RECT 119.800 6.800 120.200 7.600 ;
        RECT 121.400 7.200 121.700 7.800 ;
        RECT 123.100 7.700 124.900 7.900 ;
        RECT 123.400 7.200 123.800 7.400 ;
        RECT 125.400 7.200 125.700 7.900 ;
        RECT 121.400 6.800 121.800 7.200 ;
        RECT 122.200 7.100 122.600 7.200 ;
        RECT 123.000 7.100 123.800 7.200 ;
        RECT 122.200 6.900 123.800 7.100 ;
        RECT 122.200 6.800 123.400 6.900 ;
        RECT 124.500 6.800 125.800 7.200 ;
        RECT 126.200 6.800 126.600 7.600 ;
        RECT 120.600 5.400 121.000 6.200 ;
        RECT 121.400 5.100 121.700 6.800 ;
        RECT 123.000 6.100 123.400 6.200 ;
        RECT 123.800 6.100 124.200 6.600 ;
        RECT 123.000 5.800 124.200 6.100 ;
        RECT 124.500 5.100 124.800 6.800 ;
        RECT 126.200 6.100 126.600 6.200 ;
        RECT 127.000 6.100 127.400 7.900 ;
        RECT 128.600 7.500 129.000 9.900 ;
        RECT 130.800 9.200 131.200 9.900 ;
        RECT 130.200 8.900 131.200 9.200 ;
        RECT 133.000 8.900 133.400 9.900 ;
        RECT 135.100 9.200 135.700 9.900 ;
        RECT 135.000 8.900 135.700 9.200 ;
        RECT 130.200 8.500 130.600 8.900 ;
        RECT 133.000 8.600 133.300 8.900 ;
        RECT 131.000 8.200 131.400 8.600 ;
        RECT 131.900 8.300 133.300 8.600 ;
        RECT 135.000 8.500 135.400 8.900 ;
        RECT 131.900 8.200 132.300 8.300 ;
        RECT 129.000 7.100 129.800 7.200 ;
        RECT 131.100 7.100 131.400 8.200 ;
        RECT 135.900 7.700 136.300 7.800 ;
        RECT 137.400 7.700 137.800 9.900 ;
        RECT 138.200 7.900 138.600 9.900 ;
        RECT 140.300 9.200 140.700 9.900 ;
        RECT 140.300 8.800 141.000 9.200 ;
        RECT 140.300 8.400 140.700 8.800 ;
        RECT 140.300 7.900 141.000 8.400 ;
        RECT 135.900 7.400 137.800 7.700 ;
        RECT 138.300 7.800 138.600 7.900 ;
        RECT 138.300 7.600 139.200 7.800 ;
        RECT 138.300 7.500 140.400 7.600 ;
        RECT 133.900 7.100 134.300 7.200 ;
        RECT 137.400 7.100 137.800 7.400 ;
        RECT 138.900 7.300 140.400 7.500 ;
        RECT 140.000 7.200 140.400 7.300 ;
        RECT 138.200 7.100 138.600 7.200 ;
        RECT 129.000 6.800 134.500 7.100 ;
        RECT 130.500 6.700 130.900 6.800 ;
        RECT 126.200 5.800 127.400 6.100 ;
        RECT 129.700 6.200 130.100 6.300 ;
        RECT 129.700 5.900 132.200 6.200 ;
        RECT 131.800 5.800 132.200 5.900 ;
        RECT 125.400 5.100 125.800 5.200 ;
        RECT 120.900 4.700 121.800 5.100 ;
        RECT 124.300 4.800 124.800 5.100 ;
        RECT 125.100 4.800 125.800 5.100 ;
        RECT 120.900 1.100 121.300 4.700 ;
        RECT 124.300 1.100 124.700 4.800 ;
        RECT 125.100 4.200 125.400 4.800 ;
        RECT 125.000 3.800 125.400 4.200 ;
        RECT 127.000 1.100 127.400 5.800 ;
        RECT 128.600 5.500 131.400 5.600 ;
        RECT 128.600 5.400 131.500 5.500 ;
        RECT 128.600 5.300 133.500 5.400 ;
        RECT 127.800 4.400 128.200 5.200 ;
        RECT 128.600 1.100 129.000 5.300 ;
        RECT 131.100 5.100 133.500 5.300 ;
        RECT 130.200 4.500 132.900 4.800 ;
        RECT 130.200 4.400 130.600 4.500 ;
        RECT 132.500 4.400 132.900 4.500 ;
        RECT 133.200 4.500 133.500 5.100 ;
        RECT 134.200 5.200 134.500 6.800 ;
        RECT 137.400 6.800 138.600 7.100 ;
        RECT 139.200 6.900 139.600 7.000 ;
        RECT 135.000 6.400 135.400 6.500 ;
        RECT 135.000 6.100 136.900 6.400 ;
        RECT 136.500 6.000 136.900 6.100 ;
        RECT 135.700 5.700 136.100 5.800 ;
        RECT 137.400 5.700 137.800 6.800 ;
        RECT 138.200 6.400 138.600 6.800 ;
        RECT 139.100 6.600 139.600 6.900 ;
        RECT 139.100 6.200 139.400 6.600 ;
        RECT 139.000 5.800 139.400 6.200 ;
        RECT 135.700 5.400 137.800 5.700 ;
        RECT 140.000 5.500 140.300 7.200 ;
        RECT 140.700 6.200 141.000 7.900 ;
        RECT 141.400 7.500 141.800 9.900 ;
        RECT 143.600 9.200 144.000 9.900 ;
        RECT 143.000 8.900 144.000 9.200 ;
        RECT 145.800 8.900 146.200 9.900 ;
        RECT 147.900 9.200 148.500 9.900 ;
        RECT 147.800 8.900 148.500 9.200 ;
        RECT 143.000 8.500 143.400 8.900 ;
        RECT 145.800 8.600 146.100 8.900 ;
        RECT 143.800 7.800 144.200 8.600 ;
        RECT 144.700 8.300 146.100 8.600 ;
        RECT 147.800 8.500 148.200 8.900 ;
        RECT 144.700 8.200 145.100 8.300 ;
        RECT 141.800 7.100 142.600 7.200 ;
        RECT 143.900 7.100 144.200 7.800 ;
        RECT 148.700 7.700 149.100 7.800 ;
        RECT 150.200 7.700 150.600 9.900 ;
        RECT 148.700 7.400 150.600 7.700 ;
        RECT 146.700 7.100 147.100 7.200 ;
        RECT 141.800 6.800 147.300 7.100 ;
        RECT 143.300 6.700 143.700 6.800 ;
        RECT 140.600 5.800 141.000 6.200 ;
        RECT 142.500 6.200 142.900 6.300 ;
        RECT 142.500 5.900 145.000 6.200 ;
        RECT 144.600 5.800 145.000 5.900 ;
        RECT 134.200 4.900 135.400 5.200 ;
        RECT 133.900 4.500 134.300 4.600 ;
        RECT 133.200 4.200 134.300 4.500 ;
        RECT 135.100 4.400 135.400 4.900 ;
        RECT 135.100 4.000 135.800 4.400 ;
        RECT 131.900 3.700 132.300 3.800 ;
        RECT 133.300 3.700 133.700 3.800 ;
        RECT 130.200 3.100 130.600 3.500 ;
        RECT 131.900 3.400 133.700 3.700 ;
        RECT 133.000 3.100 133.300 3.400 ;
        RECT 135.000 3.100 135.400 3.500 ;
        RECT 130.200 2.800 131.200 3.100 ;
        RECT 130.800 1.100 131.200 2.800 ;
        RECT 133.000 1.100 133.400 3.100 ;
        RECT 135.100 1.100 135.700 3.100 ;
        RECT 137.400 1.100 137.800 5.400 ;
        RECT 139.100 5.200 140.300 5.500 ;
        RECT 139.100 3.100 139.400 5.200 ;
        RECT 140.700 5.100 141.000 5.800 ;
        RECT 139.000 1.100 139.400 3.100 ;
        RECT 140.600 1.100 141.000 5.100 ;
        RECT 141.400 5.500 144.200 5.600 ;
        RECT 141.400 5.400 144.300 5.500 ;
        RECT 141.400 5.300 146.300 5.400 ;
        RECT 141.400 1.100 141.800 5.300 ;
        RECT 143.900 5.100 146.300 5.300 ;
        RECT 143.000 4.500 145.700 4.800 ;
        RECT 143.000 4.400 143.400 4.500 ;
        RECT 145.300 4.400 145.700 4.500 ;
        RECT 146.000 4.500 146.300 5.100 ;
        RECT 147.000 5.200 147.300 6.800 ;
        RECT 147.800 6.400 148.200 6.500 ;
        RECT 147.800 6.100 149.700 6.400 ;
        RECT 149.300 6.000 149.700 6.100 ;
        RECT 148.500 5.700 148.900 5.800 ;
        RECT 150.200 5.700 150.600 7.400 ;
        RECT 148.500 5.400 150.600 5.700 ;
        RECT 147.000 4.900 148.200 5.200 ;
        RECT 146.700 4.500 147.100 4.600 ;
        RECT 146.000 4.200 147.100 4.500 ;
        RECT 147.900 4.400 148.200 4.900 ;
        RECT 147.900 4.000 148.600 4.400 ;
        RECT 150.200 4.100 150.600 5.400 ;
        RECT 152.600 7.700 153.000 9.900 ;
        RECT 154.700 9.200 155.300 9.900 ;
        RECT 154.700 8.900 155.400 9.200 ;
        RECT 157.000 8.900 157.400 9.900 ;
        RECT 159.200 9.200 159.600 9.900 ;
        RECT 159.200 8.900 160.200 9.200 ;
        RECT 155.000 8.500 155.400 8.900 ;
        RECT 157.100 8.600 157.400 8.900 ;
        RECT 157.100 8.300 158.500 8.600 ;
        RECT 158.100 8.200 158.500 8.300 ;
        RECT 159.000 7.800 159.400 8.600 ;
        RECT 159.800 8.500 160.200 8.900 ;
        RECT 154.100 7.700 154.500 7.800 ;
        RECT 152.600 7.400 154.500 7.700 ;
        RECT 152.600 5.700 153.000 7.400 ;
        RECT 156.100 7.100 156.500 7.200 ;
        RECT 159.000 7.100 159.300 7.800 ;
        RECT 161.400 7.500 161.800 9.900 ;
        RECT 163.000 8.900 163.400 9.900 ;
        RECT 162.200 7.800 162.600 8.600 ;
        RECT 163.100 7.200 163.400 8.900 ;
        RECT 164.600 7.600 165.000 9.900 ;
        RECT 164.600 7.300 165.700 7.600 ;
        RECT 160.600 7.100 161.400 7.200 ;
        RECT 155.900 6.800 161.400 7.100 ;
        RECT 163.000 6.800 163.400 7.200 ;
        RECT 155.000 6.400 155.400 6.500 ;
        RECT 153.500 6.100 155.400 6.400 ;
        RECT 153.500 6.000 153.900 6.100 ;
        RECT 154.300 5.700 154.700 5.800 ;
        RECT 152.600 5.400 154.700 5.700 ;
        RECT 152.600 4.100 153.000 5.400 ;
        RECT 155.900 5.200 156.200 6.800 ;
        RECT 159.500 6.700 159.900 6.800 ;
        RECT 160.300 6.200 160.700 6.300 ;
        RECT 158.200 5.900 160.700 6.200 ;
        RECT 158.200 5.800 158.600 5.900 ;
        RECT 159.000 5.500 161.800 5.600 ;
        RECT 158.900 5.400 161.800 5.500 ;
        RECT 155.000 4.900 156.200 5.200 ;
        RECT 156.900 5.300 161.800 5.400 ;
        RECT 156.900 5.100 159.300 5.300 ;
        RECT 155.000 4.400 155.300 4.900 ;
        RECT 150.200 3.800 153.000 4.100 ;
        RECT 154.600 4.000 155.300 4.400 ;
        RECT 156.100 4.500 156.500 4.600 ;
        RECT 156.900 4.500 157.200 5.100 ;
        RECT 156.100 4.200 157.200 4.500 ;
        RECT 157.500 4.500 160.200 4.800 ;
        RECT 157.500 4.400 157.900 4.500 ;
        RECT 159.800 4.400 160.200 4.500 ;
        RECT 144.700 3.700 145.100 3.800 ;
        RECT 146.100 3.700 146.500 3.800 ;
        RECT 143.000 3.100 143.400 3.500 ;
        RECT 144.700 3.400 146.500 3.700 ;
        RECT 145.800 3.100 146.100 3.400 ;
        RECT 147.800 3.100 148.200 3.500 ;
        RECT 143.000 2.800 144.000 3.100 ;
        RECT 143.600 1.100 144.000 2.800 ;
        RECT 145.800 1.100 146.200 3.100 ;
        RECT 147.900 1.100 148.500 3.100 ;
        RECT 150.200 1.100 150.600 3.800 ;
        RECT 152.600 1.100 153.000 3.800 ;
        RECT 156.700 3.700 157.100 3.800 ;
        RECT 158.100 3.700 158.500 3.800 ;
        RECT 155.000 3.100 155.400 3.500 ;
        RECT 156.700 3.400 158.500 3.700 ;
        RECT 157.100 3.100 157.400 3.400 ;
        RECT 159.800 3.100 160.200 3.500 ;
        RECT 154.700 1.100 155.300 3.100 ;
        RECT 157.000 1.100 157.400 3.100 ;
        RECT 159.200 2.800 160.200 3.100 ;
        RECT 159.200 1.100 159.600 2.800 ;
        RECT 161.400 1.100 161.800 5.300 ;
        RECT 163.100 5.200 163.400 6.800 ;
        RECT 163.800 5.400 164.200 6.200 ;
        RECT 165.400 5.800 165.700 7.300 ;
        RECT 166.200 6.200 166.600 9.900 ;
        RECT 167.000 8.000 167.400 9.900 ;
        RECT 168.600 8.000 169.000 9.900 ;
        RECT 167.000 7.900 169.000 8.000 ;
        RECT 169.400 8.100 169.800 9.900 ;
        RECT 171.000 8.900 171.400 9.900 ;
        RECT 170.200 8.100 170.600 8.600 ;
        RECT 171.100 8.100 171.400 8.900 ;
        RECT 167.100 7.700 168.900 7.900 ;
        RECT 169.400 7.800 170.600 8.100 ;
        RECT 171.000 7.800 172.100 8.100 ;
        RECT 167.400 7.200 167.800 7.400 ;
        RECT 169.400 7.200 169.700 7.800 ;
        RECT 171.100 7.200 171.400 7.800 ;
        RECT 167.000 6.900 167.800 7.200 ;
        RECT 167.000 6.800 167.400 6.900 ;
        RECT 168.500 6.800 169.800 7.200 ;
        RECT 171.000 6.800 171.400 7.200 ;
        RECT 171.800 7.200 172.100 7.800 ;
        RECT 172.600 7.700 173.000 9.900 ;
        RECT 174.700 9.200 175.300 9.900 ;
        RECT 174.700 8.900 175.400 9.200 ;
        RECT 177.000 8.900 177.400 9.900 ;
        RECT 179.200 9.200 179.600 9.900 ;
        RECT 179.200 8.900 180.200 9.200 ;
        RECT 175.000 8.500 175.400 8.900 ;
        RECT 177.100 8.600 177.400 8.900 ;
        RECT 177.100 8.300 178.500 8.600 ;
        RECT 178.100 8.200 178.500 8.300 ;
        RECT 179.000 8.200 179.400 8.600 ;
        RECT 179.800 8.500 180.200 8.900 ;
        RECT 174.100 7.700 174.500 7.800 ;
        RECT 172.600 7.400 174.500 7.700 ;
        RECT 171.800 6.800 172.200 7.200 ;
        RECT 165.400 5.400 166.000 5.800 ;
        RECT 163.000 5.100 163.400 5.200 ;
        RECT 165.400 5.100 165.700 5.400 ;
        RECT 166.300 5.100 166.600 6.200 ;
        RECT 167.000 6.100 167.400 6.200 ;
        RECT 167.800 6.100 168.200 6.600 ;
        RECT 167.000 5.800 168.200 6.100 ;
        RECT 168.500 5.100 168.800 6.800 ;
        RECT 169.400 5.100 169.800 5.200 ;
        RECT 171.100 5.100 171.400 6.800 ;
        RECT 171.800 5.400 172.200 6.200 ;
        RECT 172.600 5.700 173.000 7.400 ;
        RECT 176.100 7.100 176.500 7.200 ;
        RECT 179.000 7.100 179.300 8.200 ;
        RECT 181.400 7.500 181.800 9.900 ;
        RECT 183.000 8.900 183.400 9.900 ;
        RECT 182.200 8.100 182.600 8.200 ;
        RECT 183.000 8.100 183.300 8.900 ;
        RECT 182.200 7.800 183.300 8.100 ;
        RECT 183.800 7.800 184.200 8.600 ;
        RECT 183.000 7.200 183.300 7.800 ;
        RECT 184.600 7.500 185.000 9.900 ;
        RECT 186.800 9.200 187.200 9.900 ;
        RECT 186.200 8.900 187.200 9.200 ;
        RECT 189.000 8.900 189.400 9.900 ;
        RECT 191.100 9.200 191.700 9.900 ;
        RECT 191.000 8.900 191.700 9.200 ;
        RECT 193.400 9.100 193.800 9.900 ;
        RECT 194.200 9.100 194.600 9.200 ;
        RECT 186.200 8.500 186.600 8.900 ;
        RECT 189.000 8.600 189.300 8.900 ;
        RECT 187.000 8.200 187.400 8.600 ;
        RECT 187.900 8.300 189.300 8.600 ;
        RECT 191.000 8.500 191.400 8.900 ;
        RECT 193.400 8.800 194.600 9.100 ;
        RECT 187.900 8.200 188.300 8.300 ;
        RECT 180.600 7.100 181.400 7.200 ;
        RECT 175.900 6.800 181.400 7.100 ;
        RECT 183.000 6.800 183.400 7.200 ;
        RECT 185.000 7.100 185.800 7.200 ;
        RECT 187.100 7.100 187.400 8.200 ;
        RECT 191.900 7.700 192.300 7.800 ;
        RECT 193.400 7.700 193.800 8.800 ;
        RECT 191.900 7.400 193.800 7.700 ;
        RECT 189.900 7.100 190.300 7.200 ;
        RECT 185.000 6.800 190.500 7.100 ;
        RECT 175.000 6.400 175.400 6.500 ;
        RECT 173.500 6.100 175.400 6.400 ;
        RECT 175.900 6.200 176.200 6.800 ;
        RECT 179.500 6.700 179.900 6.800 ;
        RECT 180.300 6.200 180.700 6.300 ;
        RECT 173.500 6.000 173.900 6.100 ;
        RECT 175.800 5.800 176.200 6.200 ;
        RECT 178.200 5.900 180.700 6.200 ;
        RECT 178.200 5.800 178.600 5.900 ;
        RECT 174.300 5.700 174.700 5.800 ;
        RECT 172.600 5.400 174.700 5.700 ;
        RECT 163.000 4.700 163.900 5.100 ;
        RECT 163.500 1.100 163.900 4.700 ;
        RECT 164.600 4.800 165.700 5.100 ;
        RECT 164.600 1.100 165.000 4.800 ;
        RECT 166.200 1.100 166.600 5.100 ;
        RECT 168.300 4.800 168.800 5.100 ;
        RECT 169.100 4.800 169.800 5.100 ;
        RECT 168.300 1.100 168.700 4.800 ;
        RECT 169.100 4.200 169.400 4.800 ;
        RECT 171.000 4.700 171.900 5.100 ;
        RECT 169.000 3.800 169.400 4.200 ;
        RECT 171.500 1.100 171.900 4.700 ;
        RECT 172.600 1.100 173.000 5.400 ;
        RECT 175.900 5.200 176.200 5.800 ;
        RECT 179.000 5.500 181.800 5.600 ;
        RECT 178.900 5.400 181.800 5.500 ;
        RECT 182.200 5.400 182.600 6.200 ;
        RECT 175.000 4.900 176.200 5.200 ;
        RECT 176.900 5.300 181.800 5.400 ;
        RECT 176.900 5.100 179.300 5.300 ;
        RECT 175.000 4.400 175.300 4.900 ;
        RECT 174.600 4.000 175.300 4.400 ;
        RECT 176.100 4.500 176.500 4.600 ;
        RECT 176.900 4.500 177.200 5.100 ;
        RECT 176.100 4.200 177.200 4.500 ;
        RECT 177.500 4.500 180.200 4.800 ;
        RECT 177.500 4.400 177.900 4.500 ;
        RECT 179.800 4.400 180.200 4.500 ;
        RECT 176.700 3.700 177.100 3.800 ;
        RECT 178.100 3.700 178.500 3.800 ;
        RECT 175.000 3.100 175.400 3.500 ;
        RECT 176.700 3.400 178.500 3.700 ;
        RECT 177.100 3.100 177.400 3.400 ;
        RECT 179.800 3.100 180.200 3.500 ;
        RECT 174.700 1.100 175.300 3.100 ;
        RECT 177.000 1.100 177.400 3.100 ;
        RECT 179.200 2.800 180.200 3.100 ;
        RECT 179.200 1.100 179.600 2.800 ;
        RECT 181.400 1.100 181.800 5.300 ;
        RECT 183.000 5.100 183.300 6.800 ;
        RECT 186.500 6.700 186.900 6.800 ;
        RECT 185.700 6.200 186.100 6.300 ;
        RECT 185.700 5.900 188.200 6.200 ;
        RECT 187.800 5.800 188.200 5.900 ;
        RECT 184.600 5.500 187.400 5.600 ;
        RECT 184.600 5.400 187.500 5.500 ;
        RECT 184.600 5.300 189.500 5.400 ;
        RECT 182.500 4.700 183.400 5.100 ;
        RECT 182.500 1.100 182.900 4.700 ;
        RECT 184.600 1.100 185.000 5.300 ;
        RECT 187.100 5.100 189.500 5.300 ;
        RECT 186.200 4.500 188.900 4.800 ;
        RECT 186.200 4.400 186.600 4.500 ;
        RECT 188.500 4.400 188.900 4.500 ;
        RECT 189.200 4.500 189.500 5.100 ;
        RECT 190.200 5.200 190.500 6.800 ;
        RECT 191.000 6.400 191.400 6.500 ;
        RECT 191.000 6.100 192.900 6.400 ;
        RECT 192.500 6.000 192.900 6.100 ;
        RECT 191.700 5.700 192.100 5.800 ;
        RECT 193.400 5.700 193.800 7.400 ;
        RECT 191.700 5.400 193.800 5.700 ;
        RECT 190.200 4.900 191.400 5.200 ;
        RECT 189.900 4.500 190.300 4.600 ;
        RECT 189.200 4.200 190.300 4.500 ;
        RECT 191.100 4.400 191.400 4.900 ;
        RECT 191.100 4.000 191.800 4.400 ;
        RECT 187.900 3.700 188.300 3.800 ;
        RECT 189.300 3.700 189.700 3.800 ;
        RECT 186.200 3.100 186.600 3.500 ;
        RECT 187.900 3.400 189.700 3.700 ;
        RECT 189.000 3.100 189.300 3.400 ;
        RECT 191.000 3.100 191.400 3.500 ;
        RECT 186.200 2.800 187.200 3.100 ;
        RECT 186.800 1.100 187.200 2.800 ;
        RECT 189.000 1.100 189.400 3.100 ;
        RECT 191.100 1.100 191.700 3.100 ;
        RECT 193.400 1.100 193.800 5.400 ;
      LAYER via1 ;
        RECT 9.400 166.800 9.800 167.200 ;
        RECT 11.800 166.800 12.200 167.200 ;
        RECT 7.800 165.800 8.200 166.200 ;
        RECT 14.200 166.800 14.600 167.200 ;
        RECT 11.800 164.800 12.200 165.200 ;
        RECT 15.000 165.800 15.400 166.200 ;
        RECT 18.200 165.800 18.600 166.200 ;
        RECT 31.000 166.800 31.400 167.200 ;
        RECT 25.400 166.100 25.800 166.500 ;
        RECT 29.400 165.900 29.800 166.300 ;
        RECT 40.600 166.800 41.000 167.200 ;
        RECT 35.000 166.100 35.400 166.500 ;
        RECT 31.800 165.100 32.200 165.500 ;
        RECT 23.000 161.800 23.400 162.200 ;
        RECT 39.000 165.900 39.400 166.300 ;
        RECT 41.400 165.100 41.800 165.500 ;
        RECT 43.800 165.800 44.200 166.200 ;
        RECT 32.600 161.800 33.000 162.200 ;
        RECT 49.400 165.800 49.800 166.200 ;
        RECT 53.400 166.100 53.800 166.500 ;
        RECT 55.000 165.800 55.400 166.200 ;
        RECT 57.400 165.900 57.800 166.300 ;
        RECT 60.600 165.800 61.000 166.200 ;
        RECT 59.800 165.100 60.200 165.500 ;
        RECT 62.200 165.800 62.600 166.200 ;
        RECT 69.400 166.800 69.800 167.200 ;
        RECT 65.400 166.100 65.800 166.500 ;
        RECT 51.000 161.800 51.400 162.200 ;
        RECT 80.600 166.800 81.000 167.200 ;
        RECT 75.000 166.100 75.400 166.500 ;
        RECT 71.800 165.100 72.200 165.500 ;
        RECT 63.000 161.800 63.400 162.200 ;
        RECT 79.000 165.900 79.400 166.300 ;
        RECT 81.400 165.100 81.800 165.500 ;
        RECT 72.600 161.800 73.000 162.200 ;
        RECT 86.200 165.800 86.600 166.200 ;
        RECT 93.400 166.100 93.800 166.500 ;
        RECT 97.400 165.900 97.800 166.300 ;
        RECT 99.800 165.100 100.200 165.500 ;
        RECT 103.800 165.800 104.200 166.200 ;
        RECT 115.000 166.800 115.400 167.200 ;
        RECT 109.400 166.100 109.800 166.500 ;
        RECT 91.000 161.800 91.400 162.200 ;
        RECT 115.800 165.100 116.200 165.500 ;
        RECT 107.000 161.800 107.400 162.200 ;
        RECT 123.800 166.100 124.200 166.500 ;
        RECT 130.200 165.100 130.600 165.500 ;
        RECT 121.400 161.800 121.800 162.200 ;
        RECT 138.200 166.800 138.600 167.200 ;
        RECT 135.800 165.100 136.200 165.500 ;
        RECT 147.000 165.800 147.400 166.200 ;
        RECT 144.600 161.800 145.000 162.200 ;
        RECT 160.600 166.800 161.000 167.200 ;
        RECT 156.600 166.100 157.000 166.500 ;
        RECT 163.000 165.100 163.400 165.500 ;
        RECT 154.200 161.800 154.600 162.200 ;
        RECT 163.800 165.100 164.200 165.500 ;
        RECT 183.800 166.800 184.200 167.200 ;
        RECT 178.200 166.100 178.600 166.500 ;
        RECT 179.800 165.800 180.200 166.200 ;
        RECT 172.600 161.800 173.000 162.200 ;
        RECT 184.600 165.100 185.000 165.500 ;
        RECT 175.800 161.800 176.200 162.200 ;
        RECT 194.200 161.800 194.600 162.200 ;
        RECT 7.800 156.200 8.200 156.600 ;
        RECT 12.600 158.800 13.000 159.200 ;
        RECT 9.400 155.500 9.800 155.900 ;
        RECT 14.200 154.800 14.600 155.200 ;
        RECT 19.000 154.800 19.400 155.200 ;
        RECT 7.000 152.800 7.400 153.200 ;
        RECT 0.600 151.800 1.000 152.200 ;
        RECT 9.400 153.100 9.800 153.500 ;
        RECT 23.800 154.800 24.200 155.200 ;
        RECT 28.600 154.800 29.000 155.200 ;
        RECT 36.600 156.200 37.000 156.600 ;
        RECT 38.200 155.500 38.600 155.900 ;
        RECT 38.200 153.100 38.600 153.500 ;
        RECT 29.400 151.800 29.800 152.200 ;
        RECT 39.000 153.100 39.400 153.500 ;
        RECT 47.800 151.800 48.200 152.200 ;
        RECT 59.000 156.200 59.400 156.600 ;
        RECT 60.600 155.500 61.000 155.900 ;
        RECT 51.000 152.800 51.400 153.200 ;
        RECT 68.600 156.200 69.000 156.600 ;
        RECT 70.200 155.500 70.600 155.900 ;
        RECT 60.600 153.100 61.000 153.500 ;
        RECT 51.800 151.800 52.200 152.200 ;
        RECT 78.200 156.200 78.600 156.600 ;
        RECT 79.800 155.500 80.200 155.900 ;
        RECT 70.200 153.100 70.600 153.500 ;
        RECT 61.400 151.800 61.800 152.200 ;
        RECT 87.800 156.200 88.200 156.600 ;
        RECT 89.400 155.500 89.800 155.900 ;
        RECT 98.200 156.800 98.600 157.200 ;
        RECT 77.400 152.800 77.800 153.200 ;
        RECT 71.000 151.800 71.400 152.200 ;
        RECT 79.800 153.100 80.200 153.500 ;
        RECT 94.200 154.800 94.600 155.200 ;
        RECT 89.400 153.100 89.800 153.500 ;
        RECT 80.600 151.800 81.000 152.200 ;
        RECT 92.600 152.800 93.000 153.200 ;
        RECT 100.600 154.800 101.000 155.200 ;
        RECT 101.400 154.800 101.800 155.200 ;
        RECT 107.800 154.800 108.200 155.200 ;
        RECT 110.200 154.800 110.600 155.200 ;
        RECT 111.000 154.800 111.400 155.200 ;
        RECT 127.000 158.800 127.400 159.200 ;
        RECT 104.600 152.800 105.000 153.200 ;
        RECT 117.400 152.800 117.800 153.200 ;
        RECT 125.400 154.800 125.800 155.200 ;
        RECT 125.400 153.800 125.800 154.200 ;
        RECT 130.200 154.800 130.600 155.200 ;
        RECT 127.800 152.800 128.200 153.200 ;
        RECT 142.200 156.200 142.600 156.600 ;
        RECT 143.800 155.500 144.200 155.900 ;
        RECT 162.200 158.800 162.600 159.200 ;
        RECT 160.600 156.800 161.000 157.200 ;
        RECT 146.200 154.800 146.600 155.200 ;
        RECT 134.200 152.800 134.600 153.200 ;
        RECT 147.800 154.800 148.200 155.200 ;
        RECT 150.200 154.800 150.600 155.200 ;
        RECT 156.600 154.800 157.000 155.200 ;
        RECT 143.800 153.100 144.200 153.500 ;
        RECT 135.000 151.800 135.400 152.200 ;
        RECT 154.200 153.800 154.600 154.200 ;
        RECT 152.600 152.800 153.000 153.200 ;
        RECT 153.400 153.100 153.800 153.500 ;
        RECT 171.800 154.800 172.200 155.200 ;
        RECT 173.400 154.800 173.800 155.200 ;
        RECT 174.200 154.800 174.600 155.200 ;
        RECT 166.200 152.800 166.600 153.200 ;
        RECT 181.400 158.800 181.800 159.200 ;
        RECT 191.800 157.800 192.200 158.200 ;
        RECT 182.200 152.800 182.600 153.200 ;
        RECT 183.000 153.100 183.400 153.500 ;
        RECT 8.600 146.800 9.000 147.200 ;
        RECT 3.000 146.100 3.400 146.500 ;
        RECT 9.400 145.100 9.800 145.500 ;
        RECT 11.800 145.800 12.200 146.200 ;
        RECT 0.600 143.800 1.000 144.200 ;
        RECT 16.600 145.800 17.000 146.200 ;
        RECT 19.800 146.100 20.200 146.500 ;
        RECT 23.800 145.900 24.200 146.300 ;
        RECT 32.600 146.800 33.000 147.200 ;
        RECT 40.600 148.800 41.000 149.200 ;
        RECT 37.400 146.800 37.800 147.200 ;
        RECT 29.400 146.100 29.800 146.500 ;
        RECT 26.200 145.100 26.600 145.500 ;
        RECT 17.400 141.800 17.800 142.200 ;
        RECT 33.400 145.900 33.800 146.300 ;
        RECT 35.800 145.100 36.200 145.500 ;
        RECT 27.000 141.800 27.400 142.200 ;
        RECT 41.400 146.800 41.800 147.200 ;
        RECT 42.200 145.800 42.600 146.200 ;
        RECT 49.400 147.400 49.800 147.800 ;
        RECT 51.000 146.800 51.400 147.200 ;
        RECT 52.600 146.800 53.000 147.200 ;
        RECT 43.800 141.800 44.200 142.200 ;
        RECT 61.400 148.800 61.800 149.200 ;
        RECT 60.600 146.800 61.000 147.200 ;
        RECT 68.600 148.800 69.000 149.200 ;
        RECT 59.000 141.800 59.400 142.200 ;
        RECT 66.200 145.800 66.600 146.200 ;
        RECT 70.200 145.800 70.600 146.200 ;
        RECT 87.800 148.800 88.200 149.200 ;
        RECT 82.200 146.800 82.600 147.200 ;
        RECT 76.600 146.100 77.000 146.500 ;
        RECT 80.600 145.900 81.000 146.300 ;
        RECT 87.000 146.800 87.400 147.200 ;
        RECT 83.000 145.100 83.400 145.500 ;
        RECT 85.400 145.800 85.800 146.200 ;
        RECT 95.000 148.800 95.400 149.200 ;
        RECT 101.400 148.800 101.800 149.200 ;
        RECT 103.800 148.800 104.200 149.200 ;
        RECT 74.200 141.800 74.600 142.200 ;
        RECT 93.400 145.800 93.800 146.200 ;
        RECT 113.400 148.800 113.800 149.200 ;
        RECT 106.200 146.100 106.600 146.500 ;
        RECT 110.200 145.900 110.600 146.300 ;
        RECT 132.600 148.800 133.000 149.200 ;
        RECT 121.400 146.800 121.800 147.200 ;
        RECT 125.400 146.800 125.800 147.200 ;
        RECT 115.800 146.100 116.200 146.500 ;
        RECT 112.600 145.100 113.000 145.500 ;
        RECT 119.800 145.900 120.200 146.300 ;
        RECT 123.000 145.800 123.400 146.200 ;
        RECT 122.200 145.100 122.600 145.500 ;
        RECT 113.400 141.800 113.800 142.200 ;
        RECT 147.800 148.800 148.200 149.200 ;
        RECT 159.800 148.800 160.200 149.200 ;
        RECT 135.000 146.100 135.400 146.500 ;
        RECT 139.000 145.900 139.400 146.300 ;
        RECT 151.800 146.800 152.200 147.200 ;
        RECT 162.200 148.800 162.600 149.200 ;
        RECT 141.400 145.100 141.800 145.500 ;
        RECT 132.600 141.800 133.000 142.200 ;
        RECT 151.000 145.100 151.400 145.500 ;
        RECT 175.800 146.800 176.200 147.200 ;
        RECT 162.200 144.800 162.600 145.200 ;
        RECT 161.400 141.800 161.800 142.200 ;
        RECT 165.400 144.800 165.800 145.200 ;
        RECT 170.200 145.800 170.600 146.200 ;
        RECT 175.000 145.900 175.400 146.300 ;
        RECT 171.000 144.800 171.400 145.200 ;
        RECT 172.600 145.100 173.000 145.500 ;
        RECT 183.000 146.800 183.400 147.200 ;
        RECT 184.600 145.900 185.000 146.300 ;
        RECT 181.400 142.800 181.800 143.200 ;
        RECT 182.200 145.100 182.600 145.500 ;
        RECT 191.000 142.800 191.400 143.200 ;
        RECT 0.600 136.800 1.000 137.200 ;
        RECT 7.800 136.200 8.200 136.600 ;
        RECT 9.400 135.500 9.800 135.900 ;
        RECT 19.000 136.800 19.400 137.200 ;
        RECT 13.400 134.800 13.800 135.200 ;
        RECT 9.400 133.100 9.800 133.500 ;
        RECT 10.200 133.100 10.600 133.500 ;
        RECT 22.200 134.800 22.600 135.200 ;
        RECT 23.000 134.800 23.400 135.200 ;
        RECT 26.200 134.800 26.600 135.200 ;
        RECT 19.800 132.800 20.200 133.200 ;
        RECT 44.600 136.800 45.000 137.200 ;
        RECT 51.000 138.800 51.400 139.200 ;
        RECT 35.000 134.800 35.400 135.200 ;
        RECT 35.800 134.800 36.200 135.200 ;
        RECT 43.000 135.800 43.400 136.200 ;
        RECT 48.600 135.900 49.000 136.300 ;
        RECT 54.200 138.800 54.600 139.200 ;
        RECT 61.400 138.800 61.800 139.200 ;
        RECT 67.000 138.800 67.400 139.200 ;
        RECT 64.600 136.800 65.000 137.200 ;
        RECT 67.800 136.800 68.200 137.200 ;
        RECT 38.200 134.800 38.600 135.200 ;
        RECT 37.400 133.800 37.800 134.200 ;
        RECT 31.000 132.800 31.400 133.200 ;
        RECT 30.200 131.800 30.600 132.200 ;
        RECT 39.000 133.800 39.400 134.200 ;
        RECT 44.600 134.800 45.000 135.200 ;
        RECT 40.600 131.800 41.000 132.200 ;
        RECT 48.600 133.100 49.000 133.500 ;
        RECT 52.600 133.800 53.000 134.200 ;
        RECT 51.000 133.200 51.400 133.600 ;
        RECT 55.800 134.800 56.200 135.200 ;
        RECT 57.400 134.800 57.800 135.200 ;
        RECT 63.000 135.800 63.400 136.200 ;
        RECT 66.200 135.800 66.600 136.200 ;
        RECT 61.400 134.800 61.800 135.200 ;
        RECT 62.200 133.800 62.600 134.200 ;
        RECT 69.400 133.800 69.800 134.200 ;
        RECT 73.400 136.800 73.800 137.200 ;
        RECT 78.200 138.800 78.600 139.200 ;
        RECT 71.800 135.800 72.200 136.200 ;
        RECT 75.700 135.900 76.100 136.300 ;
        RECT 83.000 138.800 83.400 139.200 ;
        RECT 80.600 134.800 81.000 135.200 ;
        RECT 74.200 133.800 74.600 134.200 ;
        RECT 75.700 133.100 76.100 133.500 ;
        RECT 81.400 134.800 81.800 135.200 ;
        RECT 79.800 133.800 80.200 134.200 ;
        RECT 94.200 138.800 94.600 139.200 ;
        RECT 90.200 134.800 90.600 135.200 ;
        RECT 103.800 138.800 104.200 139.200 ;
        RECT 108.600 138.800 109.000 139.200 ;
        RECT 91.000 133.800 91.400 134.200 ;
        RECT 96.600 134.800 97.000 135.200 ;
        RECT 87.000 131.800 87.400 132.200 ;
        RECT 100.600 134.800 101.000 135.200 ;
        RECT 101.400 134.800 101.800 135.200 ;
        RECT 111.000 134.800 111.400 135.200 ;
        RECT 111.000 132.800 111.400 133.200 ;
        RECT 115.000 138.800 115.400 139.200 ;
        RECT 119.800 138.800 120.200 139.200 ;
        RECT 117.400 134.800 117.800 135.200 ;
        RECT 129.400 138.800 129.800 139.200 ;
        RECT 131.800 136.800 132.200 137.200 ;
        RECT 125.400 134.800 125.800 135.200 ;
        RECT 126.200 134.800 126.600 135.200 ;
        RECT 127.000 134.800 127.400 135.200 ;
        RECT 127.800 134.800 128.200 135.200 ;
        RECT 131.000 134.800 131.400 135.200 ;
        RECT 135.800 134.800 136.200 135.200 ;
        RECT 137.400 133.800 137.800 134.200 ;
        RECT 139.800 133.800 140.200 134.200 ;
        RECT 140.600 132.800 141.000 133.200 ;
        RECT 143.000 133.800 143.400 134.200 ;
        RECT 143.800 133.800 144.200 134.200 ;
        RECT 147.800 134.800 148.200 135.200 ;
        RECT 153.400 134.800 153.800 135.200 ;
        RECT 155.800 133.800 156.200 134.200 ;
        RECT 142.200 131.800 142.600 132.200 ;
        RECT 155.000 131.800 155.400 132.200 ;
        RECT 156.600 131.800 157.000 132.200 ;
        RECT 161.400 134.800 161.800 135.200 ;
        RECT 163.800 135.800 164.200 136.200 ;
        RECT 165.400 134.800 165.800 135.200 ;
        RECT 162.200 133.800 162.600 134.200 ;
        RECT 164.600 133.800 165.000 134.200 ;
        RECT 166.200 133.800 166.600 134.200 ;
        RECT 159.000 131.800 159.400 132.200 ;
        RECT 170.200 133.100 170.600 133.500 ;
        RECT 187.000 136.200 187.400 136.600 ;
        RECT 188.600 135.500 189.000 135.900 ;
        RECT 191.800 134.800 192.200 135.200 ;
        RECT 188.600 133.100 189.000 133.500 ;
        RECT 8.600 126.800 9.000 127.200 ;
        RECT 3.000 126.100 3.400 126.500 ;
        RECT 14.200 126.800 14.600 127.200 ;
        RECT 28.600 128.800 29.000 129.200 ;
        RECT 18.200 126.800 18.600 127.200 ;
        RECT 30.200 128.800 30.600 129.200 ;
        RECT 12.600 126.100 13.000 126.500 ;
        RECT 9.400 125.100 9.800 125.500 ;
        RECT 0.600 123.800 1.000 124.200 ;
        RECT 16.600 125.900 17.000 126.300 ;
        RECT 23.800 125.800 24.200 126.200 ;
        RECT 19.000 125.100 19.400 125.500 ;
        RECT 10.200 121.800 10.600 122.200 ;
        RECT 19.800 125.100 20.200 125.500 ;
        RECT 28.600 121.800 29.000 122.200 ;
        RECT 32.600 125.800 33.000 126.200 ;
        RECT 33.400 124.800 33.800 125.200 ;
        RECT 37.400 125.800 37.800 126.200 ;
        RECT 39.800 125.800 40.200 126.200 ;
        RECT 42.200 125.800 42.600 126.200 ;
        RECT 50.200 125.800 50.600 126.200 ;
        RECT 65.400 128.800 65.800 129.200 ;
        RECT 39.800 123.800 40.200 124.200 ;
        RECT 36.600 121.800 37.000 122.200 ;
        RECT 42.200 122.800 42.600 123.200 ;
        RECT 59.800 124.800 60.200 125.200 ;
        RECT 55.000 121.800 55.400 122.200 ;
        RECT 72.600 127.800 73.000 128.200 ;
        RECT 66.200 125.800 66.600 126.200 ;
        RECT 67.800 125.800 68.200 126.200 ;
        RECT 63.000 124.800 63.400 125.200 ;
        RECT 79.800 125.800 80.200 126.200 ;
        RECT 82.200 124.800 82.600 125.200 ;
        RECT 103.000 128.800 103.400 129.200 ;
        RECT 110.200 128.800 110.600 129.200 ;
        RECT 99.000 126.800 99.400 127.200 ;
        RECT 93.400 126.100 93.800 126.500 ;
        RECT 99.800 125.100 100.200 125.500 ;
        RECT 91.000 122.800 91.400 123.200 ;
        RECT 111.800 125.800 112.200 126.200 ;
        RECT 115.800 125.800 116.200 126.200 ;
        RECT 115.000 121.800 115.400 122.200 ;
        RECT 119.800 127.800 120.200 128.200 ;
        RECT 122.200 125.800 122.600 126.200 ;
        RECT 134.200 128.800 134.600 129.200 ;
        RECT 127.800 121.800 128.200 122.200 ;
        RECT 131.000 121.800 131.400 122.200 ;
        RECT 142.200 126.800 142.600 127.200 ;
        RECT 141.400 125.800 141.800 126.200 ;
        RECT 139.800 124.800 140.200 125.200 ;
        RECT 143.000 125.800 143.400 126.200 ;
        RECT 145.400 125.800 145.800 126.200 ;
        RECT 145.400 124.800 145.800 125.200 ;
        RECT 147.800 125.800 148.200 126.200 ;
        RECT 150.200 125.800 150.600 126.200 ;
        RECT 157.400 125.800 157.800 126.200 ;
        RECT 161.400 125.800 161.800 126.200 ;
        RECT 170.200 127.400 170.600 127.800 ;
        RECT 171.800 126.800 172.200 127.200 ;
        RECT 184.600 127.800 185.000 128.200 ;
        RECT 175.000 126.100 175.400 126.500 ;
        RECT 183.000 125.800 183.400 126.200 ;
        RECT 181.400 125.100 181.800 125.500 ;
        RECT 172.600 121.800 173.000 122.200 ;
        RECT 190.200 125.800 190.600 126.200 ;
        RECT 195.000 125.800 195.400 126.200 ;
        RECT 195.000 121.800 195.400 122.200 ;
        RECT 0.600 118.800 1.000 119.200 ;
        RECT 7.800 116.200 8.200 116.600 ;
        RECT 9.400 115.500 9.800 115.900 ;
        RECT 9.400 113.100 9.800 113.500 ;
        RECT 10.200 112.800 10.600 113.200 ;
        RECT 19.000 114.800 19.400 115.200 ;
        RECT 11.000 111.800 11.400 112.200 ;
        RECT 15.800 113.100 16.200 113.500 ;
        RECT 15.000 111.800 15.400 112.200 ;
        RECT 18.200 112.800 18.600 113.200 ;
        RECT 32.600 116.200 33.000 116.600 ;
        RECT 34.200 115.500 34.600 115.900 ;
        RECT 35.800 114.800 36.200 115.200 ;
        RECT 43.800 118.800 44.200 119.200 ;
        RECT 43.000 116.800 43.400 117.200 ;
        RECT 44.600 116.800 45.000 117.200 ;
        RECT 49.400 116.800 49.800 117.200 ;
        RECT 51.000 116.800 51.400 117.200 ;
        RECT 52.600 116.800 53.000 117.200 ;
        RECT 34.200 113.100 34.600 113.500 ;
        RECT 47.800 115.800 48.200 116.200 ;
        RECT 45.400 114.800 45.800 115.200 ;
        RECT 51.000 115.800 51.400 116.200 ;
        RECT 50.200 114.800 50.600 115.200 ;
        RECT 54.200 115.800 54.600 116.200 ;
        RECT 55.800 115.800 56.200 116.200 ;
        RECT 53.400 114.800 53.800 115.200 ;
        RECT 25.400 111.800 25.800 112.200 ;
        RECT 39.000 112.800 39.400 113.200 ;
        RECT 41.400 112.800 41.800 113.200 ;
        RECT 63.000 115.800 63.400 116.200 ;
        RECT 60.600 114.800 61.000 115.200 ;
        RECT 58.200 113.800 58.600 114.200 ;
        RECT 57.400 112.800 57.800 113.200 ;
        RECT 61.400 113.800 61.800 114.200 ;
        RECT 69.400 118.800 69.800 119.200 ;
        RECT 63.000 112.800 63.400 113.200 ;
        RECT 67.000 112.800 67.400 113.200 ;
        RECT 76.600 116.200 77.000 116.600 ;
        RECT 78.200 115.500 78.600 115.900 ;
        RECT 81.400 114.800 81.800 115.200 ;
        RECT 78.200 113.100 78.600 113.500 ;
        RECT 67.800 111.800 68.200 112.200 ;
        RECT 79.800 112.800 80.200 113.200 ;
        RECT 86.200 114.800 86.600 115.200 ;
        RECT 87.000 114.800 87.400 115.200 ;
        RECT 85.400 113.800 85.800 114.200 ;
        RECT 102.200 116.200 102.600 116.600 ;
        RECT 103.800 115.500 104.200 115.900 ;
        RECT 107.800 114.800 108.200 115.200 ;
        RECT 92.600 112.800 93.000 113.200 ;
        RECT 103.800 113.100 104.200 113.500 ;
        RECT 91.800 111.800 92.200 112.200 ;
        RECT 95.000 111.800 95.400 112.200 ;
        RECT 104.600 113.100 105.000 113.500 ;
        RECT 114.200 116.800 114.600 117.200 ;
        RECT 121.400 116.200 121.800 116.600 ;
        RECT 123.000 115.500 123.400 115.900 ;
        RECT 127.800 115.800 128.200 116.200 ;
        RECT 125.400 113.800 125.800 114.200 ;
        RECT 129.400 114.800 129.800 115.200 ;
        RECT 130.200 114.800 130.600 115.200 ;
        RECT 123.000 113.100 123.400 113.500 ;
        RECT 123.800 112.800 124.200 113.200 ;
        RECT 133.400 112.800 133.800 113.200 ;
        RECT 131.800 111.800 132.200 112.200 ;
        RECT 135.800 113.800 136.200 114.200 ;
        RECT 139.800 114.800 140.200 115.200 ;
        RECT 143.000 118.800 143.400 119.200 ;
        RECT 142.200 112.800 142.600 113.200 ;
        RECT 153.400 116.200 153.800 116.600 ;
        RECT 155.000 115.500 155.400 115.900 ;
        RECT 145.400 112.800 145.800 113.200 ;
        RECT 155.000 113.100 155.400 113.500 ;
        RECT 146.200 111.800 146.600 112.200 ;
        RECT 166.200 116.200 166.600 116.600 ;
        RECT 167.800 115.500 168.200 115.900 ;
        RECT 168.600 116.800 169.000 117.200 ;
        RECT 175.800 116.200 176.200 116.600 ;
        RECT 177.400 115.500 177.800 115.900 ;
        RECT 179.800 115.800 180.200 116.200 ;
        RECT 167.800 113.100 168.200 113.500 ;
        RECT 158.200 111.800 158.600 112.200 ;
        RECT 159.000 111.800 159.400 112.200 ;
        RECT 182.200 114.800 182.600 115.200 ;
        RECT 184.600 114.800 185.000 115.200 ;
        RECT 186.200 114.800 186.600 115.200 ;
        RECT 177.400 113.100 177.800 113.500 ;
        RECT 185.400 113.800 185.800 114.200 ;
        RECT 2.200 104.800 2.600 105.200 ;
        RECT 5.400 105.800 5.800 106.200 ;
        RECT 7.800 106.800 8.200 107.200 ;
        RECT 11.000 105.800 11.400 106.200 ;
        RECT 13.400 106.800 13.800 107.200 ;
        RECT 12.600 105.800 13.000 106.200 ;
        RECT 12.600 103.800 13.000 104.200 ;
        RECT 15.800 101.800 16.200 102.200 ;
        RECT 19.000 104.800 19.400 105.200 ;
        RECT 22.200 105.800 22.600 106.200 ;
        RECT 29.400 106.800 29.800 107.200 ;
        RECT 27.000 101.800 27.400 102.200 ;
        RECT 31.800 104.800 32.200 105.200 ;
        RECT 44.600 107.800 45.000 108.200 ;
        RECT 39.000 104.800 39.400 105.200 ;
        RECT 53.400 105.800 53.800 106.200 ;
        RECT 40.600 102.800 41.000 103.200 ;
        RECT 51.800 101.800 52.200 102.200 ;
        RECT 57.400 105.800 57.800 106.200 ;
        RECT 70.200 108.800 70.600 109.200 ;
        RECT 64.600 106.800 65.000 107.200 ;
        RECT 60.600 104.800 61.000 105.200 ;
        RECT 67.800 106.800 68.200 107.200 ;
        RECT 67.000 105.800 67.400 106.200 ;
        RECT 76.600 108.800 77.000 109.200 ;
        RECT 73.400 105.800 73.800 106.200 ;
        RECT 83.000 108.800 83.400 109.200 ;
        RECT 94.200 108.800 94.600 109.200 ;
        RECT 91.000 106.800 91.400 107.200 ;
        RECT 85.400 106.100 85.800 106.500 ;
        RECT 89.400 105.900 89.800 106.300 ;
        RECT 99.000 106.800 99.400 107.200 ;
        RECT 103.800 108.800 104.200 109.200 ;
        RECT 102.200 106.800 102.600 107.200 ;
        RECT 96.600 106.100 97.000 106.500 ;
        RECT 91.800 105.100 92.200 105.500 ;
        RECT 116.600 108.800 117.000 109.200 ;
        RECT 106.200 106.100 106.600 106.500 ;
        RECT 110.200 105.900 110.600 106.300 ;
        RECT 136.600 108.800 137.000 109.200 ;
        RECT 103.000 105.100 103.400 105.500 ;
        RECT 112.600 105.100 113.000 105.500 ;
        RECT 115.000 105.800 115.400 106.200 ;
        RECT 128.600 106.800 129.000 107.200 ;
        RECT 146.200 108.800 146.600 109.200 ;
        RECT 126.200 105.800 126.600 106.200 ;
        RECT 127.800 105.100 128.200 105.500 ;
        RECT 125.400 101.800 125.800 102.200 ;
        RECT 138.200 106.800 138.600 107.200 ;
        RECT 141.400 105.800 141.800 106.200 ;
        RECT 137.400 105.100 137.800 105.500 ;
        RECT 149.400 104.800 149.800 105.200 ;
        RECT 158.200 106.800 158.600 107.200 ;
        RECT 157.400 105.800 157.800 106.200 ;
        RECT 163.800 105.800 164.200 106.200 ;
        RECT 167.000 106.800 167.400 107.200 ;
        RECT 180.600 108.800 181.000 109.200 ;
        RECT 184.600 108.800 185.000 109.200 ;
        RECT 171.800 105.800 172.200 106.200 ;
        RECT 189.400 108.800 189.800 109.200 ;
        RECT 183.000 105.800 183.400 106.200 ;
        RECT 187.000 105.800 187.400 106.200 ;
        RECT 180.600 101.800 181.000 102.200 ;
        RECT 190.200 105.800 190.600 106.200 ;
        RECT 3.000 94.800 3.400 95.200 ;
        RECT 5.400 94.800 5.800 95.200 ;
        RECT 8.700 95.900 9.100 96.300 ;
        RECT 13.400 98.800 13.800 99.200 ;
        RECT 9.300 94.900 9.700 95.300 ;
        RECT 7.000 92.800 7.400 93.200 ;
        RECT 8.700 93.100 9.100 93.500 ;
        RECT 12.600 93.800 13.000 94.200 ;
        RECT 20.600 96.200 21.000 96.600 ;
        RECT 22.200 95.500 22.600 95.900 ;
        RECT 26.200 94.800 26.600 95.200 ;
        RECT 11.000 91.800 11.400 92.200 ;
        RECT 25.400 93.800 25.800 94.200 ;
        RECT 27.000 93.800 27.400 94.200 ;
        RECT 22.200 93.100 22.600 93.500 ;
        RECT 33.400 94.800 33.800 95.200 ;
        RECT 36.600 94.800 37.000 95.200 ;
        RECT 34.200 93.800 34.600 94.200 ;
        RECT 49.400 95.900 49.800 96.300 ;
        RECT 43.800 93.800 44.200 94.200 ;
        RECT 46.200 93.800 46.600 94.200 ;
        RECT 44.600 91.800 45.000 92.200 ;
        RECT 49.400 93.100 49.800 93.500 ;
        RECT 53.400 93.800 53.800 94.200 ;
        RECT 51.800 93.200 52.200 93.600 ;
        RECT 63.800 95.900 64.200 96.300 ;
        RECT 55.800 93.800 56.200 94.200 ;
        RECT 58.200 92.800 58.600 93.200 ;
        RECT 63.800 93.100 64.200 93.500 ;
        RECT 67.800 93.800 68.200 94.200 ;
        RECT 71.000 94.800 71.400 95.200 ;
        RECT 73.400 94.800 73.800 95.200 ;
        RECT 74.200 94.800 74.600 95.200 ;
        RECT 77.400 94.800 77.800 95.200 ;
        RECT 66.200 93.200 66.600 93.600 ;
        RECT 68.600 92.800 69.000 93.200 ;
        RECT 80.600 94.800 81.000 95.200 ;
        RECT 81.400 94.800 81.800 95.200 ;
        RECT 87.800 97.800 88.200 98.200 ;
        RECT 79.800 92.800 80.200 93.200 ;
        RECT 79.000 91.800 79.400 92.200 ;
        RECT 95.000 96.200 95.400 96.600 ;
        RECT 96.600 95.500 97.000 95.900 ;
        RECT 104.600 98.800 105.000 99.200 ;
        RECT 87.000 92.800 87.400 93.200 ;
        RECT 108.600 94.800 109.000 95.200 ;
        RECT 109.400 94.800 109.800 95.200 ;
        RECT 96.600 93.100 97.000 93.500 ;
        RECT 87.800 91.800 88.200 92.200 ;
        RECT 106.200 92.800 106.600 93.200 ;
        RECT 104.600 91.800 105.000 92.200 ;
        RECT 107.000 91.800 107.400 92.200 ;
        RECT 115.800 93.800 116.200 94.200 ;
        RECT 119.000 97.800 119.400 98.200 ;
        RECT 118.200 93.800 118.600 94.200 ;
        RECT 122.200 94.800 122.600 95.200 ;
        RECT 126.200 95.900 126.600 96.300 ;
        RECT 138.300 95.900 138.700 96.300 ;
        RECT 143.000 98.800 143.400 99.200 ;
        RECT 119.800 92.800 120.200 93.200 ;
        RECT 124.600 92.800 125.000 93.200 ;
        RECT 126.200 93.100 126.600 93.500 ;
        RECT 130.200 93.800 130.600 94.200 ;
        RECT 133.400 93.800 133.800 94.200 ;
        RECT 128.600 93.200 129.000 93.600 ;
        RECT 128.600 91.800 129.000 92.200 ;
        RECT 138.900 94.900 139.300 95.300 ;
        RECT 138.300 93.100 138.700 93.500 ;
        RECT 142.200 93.800 142.600 94.200 ;
        RECT 150.200 96.200 150.600 96.600 ;
        RECT 151.800 95.500 152.200 95.900 ;
        RECT 154.200 98.800 154.600 99.200 ;
        RECT 143.000 92.800 143.400 93.200 ;
        RECT 161.400 96.200 161.800 96.600 ;
        RECT 163.000 95.500 163.400 95.900 ;
        RECT 172.600 96.800 173.000 97.200 ;
        RECT 151.800 93.100 152.200 93.500 ;
        RECT 163.000 93.100 163.400 93.500 ;
        RECT 163.800 93.100 164.200 93.500 ;
        RECT 180.600 96.200 181.000 96.600 ;
        RECT 182.200 95.500 182.600 95.900 ;
        RECT 183.800 93.800 184.200 94.200 ;
        RECT 182.200 93.100 182.600 93.500 ;
        RECT 173.400 91.800 173.800 92.200 ;
        RECT 183.000 93.100 183.400 93.500 ;
        RECT 191.800 91.800 192.200 92.200 ;
        RECT 12.600 88.800 13.000 89.200 ;
        RECT 3.800 85.800 4.200 86.200 ;
        RECT 2.200 84.800 2.600 85.200 ;
        RECT 7.800 85.800 8.200 86.200 ;
        RECT 5.400 81.800 5.800 82.200 ;
        RECT 11.800 85.800 12.200 86.200 ;
        RECT 18.200 86.800 18.600 87.200 ;
        RECT 23.000 88.800 23.400 89.200 ;
        RECT 27.000 88.800 27.400 89.200 ;
        RECT 15.000 86.100 15.400 86.500 ;
        RECT 10.200 81.800 10.600 82.200 ;
        RECT 19.000 85.900 19.400 86.300 ;
        RECT 21.400 85.100 21.800 85.500 ;
        RECT 25.400 85.800 25.800 86.200 ;
        RECT 34.200 88.800 34.600 89.200 ;
        RECT 34.200 84.800 34.600 85.200 ;
        RECT 38.200 84.800 38.600 85.200 ;
        RECT 51.800 88.800 52.200 89.200 ;
        RECT 40.600 84.800 41.000 85.200 ;
        RECT 53.400 86.800 53.800 87.200 ;
        RECT 62.200 88.800 62.600 89.200 ;
        RECT 46.200 85.800 46.600 86.200 ;
        RECT 43.000 83.800 43.400 84.200 ;
        RECT 56.600 85.800 57.000 86.200 ;
        RECT 72.600 88.800 73.000 89.200 ;
        RECT 74.200 88.800 74.600 89.200 ;
        RECT 70.200 86.800 70.600 87.200 ;
        RECT 64.600 86.100 65.000 86.500 ;
        RECT 61.400 81.800 61.800 82.200 ;
        RECT 68.600 85.900 69.000 86.300 ;
        RECT 71.000 85.100 71.400 85.500 ;
        RECT 71.800 84.800 72.200 85.200 ;
        RECT 84.600 88.800 85.000 89.200 ;
        RECT 87.000 88.800 87.400 89.200 ;
        RECT 82.200 86.800 82.600 87.200 ;
        RECT 76.600 86.100 77.000 86.500 ;
        RECT 83.000 85.100 83.400 85.500 ;
        RECT 86.200 85.800 86.600 86.200 ;
        RECT 95.000 86.800 95.400 87.200 ;
        RECT 89.400 86.100 89.800 86.500 ;
        RECT 93.400 85.900 93.800 86.300 ;
        RECT 106.200 86.800 106.600 87.200 ;
        RECT 100.600 86.100 101.000 86.500 ;
        RECT 95.800 85.100 96.200 85.500 ;
        RECT 104.600 85.900 105.000 86.300 ;
        RECT 120.600 88.800 121.000 89.200 ;
        RECT 110.200 86.100 110.600 86.500 ;
        RECT 107.000 85.100 107.400 85.500 ;
        RECT 98.200 81.800 98.600 82.200 ;
        RECT 116.600 85.100 117.000 85.500 ;
        RECT 119.000 85.800 119.400 86.200 ;
        RECT 107.800 81.800 108.200 82.200 ;
        RECT 119.800 84.800 120.200 85.200 ;
        RECT 119.000 81.800 119.400 82.200 ;
        RECT 127.000 88.800 127.400 89.200 ;
        RECT 125.400 85.800 125.800 86.200 ;
        RECT 133.400 86.800 133.800 87.200 ;
        RECT 135.000 86.800 135.400 87.200 ;
        RECT 138.200 86.800 138.600 87.200 ;
        RECT 145.400 88.800 145.800 89.200 ;
        RECT 129.400 86.100 129.800 86.500 ;
        RECT 135.800 85.100 136.200 85.500 ;
        RECT 138.200 85.800 138.600 86.200 ;
        RECT 151.000 86.800 151.400 87.200 ;
        RECT 147.800 86.100 148.200 86.500 ;
        RECT 140.600 84.800 141.000 85.200 ;
        RECT 159.800 88.800 160.200 89.200 ;
        RECT 154.200 85.100 154.600 85.500 ;
        RECT 164.600 85.800 165.000 86.200 ;
        RECT 166.200 85.800 166.600 86.200 ;
        RECT 167.800 85.800 168.200 86.200 ;
        RECT 174.200 85.800 174.600 86.200 ;
        RECT 164.600 81.800 165.000 82.200 ;
        RECT 167.000 81.800 167.400 82.200 ;
        RECT 175.800 84.800 176.200 85.200 ;
        RECT 178.200 85.800 178.600 86.200 ;
        RECT 179.000 85.800 179.400 86.200 ;
        RECT 184.600 87.400 185.000 87.800 ;
        RECT 186.200 86.800 186.600 87.200 ;
        RECT 178.200 81.800 178.600 82.200 ;
        RECT 10.200 78.800 10.600 79.200 ;
        RECT 7.800 73.800 8.200 74.200 ;
        RECT 17.400 76.200 17.800 76.600 ;
        RECT 19.000 75.500 19.400 75.900 ;
        RECT 28.600 78.800 29.000 79.200 ;
        RECT 23.000 74.800 23.400 75.200 ;
        RECT 31.800 78.800 32.200 79.200 ;
        RECT 9.400 72.800 9.800 73.200 ;
        RECT 19.000 73.100 19.400 73.500 ;
        RECT 10.200 71.800 10.600 72.200 ;
        RECT 19.800 73.100 20.200 73.500 ;
        RECT 29.400 72.800 29.800 73.200 ;
        RECT 30.200 71.800 30.600 72.200 ;
        RECT 39.000 76.200 39.400 76.600 ;
        RECT 40.600 75.500 41.000 75.900 ;
        RECT 40.600 73.100 41.000 73.500 ;
        RECT 31.800 71.800 32.200 72.200 ;
        RECT 41.400 72.800 41.800 73.200 ;
        RECT 43.800 73.800 44.200 74.200 ;
        RECT 49.400 74.800 49.800 75.200 ;
        RECT 47.000 72.800 47.400 73.200 ;
        RECT 49.400 72.800 49.800 73.200 ;
        RECT 51.000 72.800 51.400 73.200 ;
        RECT 55.800 75.800 56.200 76.200 ;
        RECT 59.800 78.800 60.200 79.200 ;
        RECT 64.600 76.800 65.000 77.200 ;
        RECT 55.800 74.800 56.200 75.200 ;
        RECT 53.400 73.800 53.800 74.200 ;
        RECT 56.600 73.800 57.000 74.200 ;
        RECT 52.600 71.800 53.000 72.200 ;
        RECT 59.800 71.800 60.200 72.200 ;
        RECT 66.200 75.800 66.600 76.200 ;
        RECT 65.400 74.800 65.800 75.200 ;
        RECT 62.200 71.800 62.600 72.200 ;
        RECT 74.200 76.200 74.600 76.600 ;
        RECT 75.800 75.500 76.200 75.900 ;
        RECT 83.000 75.800 83.400 76.200 ;
        RECT 75.800 73.100 76.200 73.500 ;
        RECT 67.000 71.800 67.400 72.200 ;
        RECT 80.600 74.800 81.000 75.200 ;
        RECT 84.600 74.800 85.000 75.200 ;
        RECT 87.800 74.800 88.200 75.200 ;
        RECT 78.200 72.800 78.600 73.200 ;
        RECT 85.400 73.800 85.800 74.200 ;
        RECT 83.000 72.800 83.400 73.200 ;
        RECT 91.800 74.800 92.200 75.200 ;
        RECT 100.600 78.800 101.000 79.200 ;
        RECT 103.000 78.800 103.400 79.200 ;
        RECT 95.800 74.800 96.200 75.200 ;
        RECT 96.600 74.800 97.000 75.200 ;
        RECT 86.200 71.800 86.600 72.200 ;
        RECT 115.000 78.800 115.400 79.200 ;
        RECT 109.400 74.800 109.800 75.200 ;
        RECT 123.000 75.800 123.400 76.200 ;
        RECT 105.400 73.800 105.800 74.200 ;
        RECT 106.200 73.100 106.600 73.500 ;
        RECT 119.000 74.800 119.400 75.200 ;
        RECT 115.800 73.100 116.200 73.500 ;
        RECT 137.400 78.800 137.800 79.200 ;
        RECT 135.000 73.800 135.400 74.200 ;
        RECT 142.200 74.800 142.600 75.200 ;
        RECT 124.600 71.800 125.000 72.200 ;
        RECT 127.000 72.800 127.400 73.200 ;
        RECT 139.000 73.100 139.400 73.500 ;
        RECT 147.800 71.800 148.200 72.200 ;
        RECT 153.400 78.800 153.800 79.200 ;
        RECT 152.600 72.800 153.000 73.200 ;
        RECT 163.000 78.800 163.400 79.200 ;
        RECT 158.200 74.800 158.600 75.200 ;
        RECT 155.000 73.800 155.400 74.200 ;
        RECT 154.200 73.100 154.600 73.500 ;
        RECT 165.400 74.800 165.800 75.200 ;
        RECT 163.000 72.800 163.400 73.200 ;
        RECT 166.200 73.800 166.600 74.200 ;
        RECT 165.400 72.800 165.800 73.200 ;
        RECT 168.600 72.800 169.000 73.200 ;
        RECT 172.600 73.800 173.000 74.200 ;
        RECT 173.400 72.800 173.800 73.200 ;
        RECT 176.600 72.800 177.000 73.200 ;
        RECT 185.400 73.800 185.800 74.200 ;
        RECT 175.800 71.800 176.200 72.200 ;
        RECT 178.200 71.800 178.600 72.200 ;
        RECT 183.800 72.800 184.200 73.200 ;
        RECT 184.600 73.100 185.000 73.500 ;
        RECT 193.400 71.800 193.800 72.200 ;
        RECT 10.200 68.800 10.600 69.200 ;
        RECT 9.400 66.800 9.800 67.200 ;
        RECT 18.200 66.800 18.600 67.200 ;
        RECT 33.400 68.800 33.800 69.200 ;
        RECT 27.000 66.800 27.400 67.200 ;
        RECT 12.600 66.100 13.000 66.500 ;
        RECT 8.600 61.800 9.000 62.200 ;
        RECT 16.600 65.900 17.000 66.300 ;
        RECT 19.000 65.100 19.400 65.500 ;
        RECT 22.200 65.800 22.600 66.200 ;
        RECT 29.400 65.800 29.800 66.200 ;
        RECT 24.600 65.100 25.000 65.500 ;
        RECT 48.600 68.800 49.000 69.200 ;
        RECT 39.800 66.800 40.200 67.200 ;
        RECT 36.600 65.800 37.000 66.200 ;
        RECT 39.000 65.100 39.400 65.500 ;
        RECT 48.600 61.800 49.000 62.200 ;
        RECT 55.000 66.800 55.400 67.200 ;
        RECT 63.000 68.800 63.400 69.200 ;
        RECT 60.600 65.800 61.000 66.200 ;
        RECT 77.400 68.800 77.800 69.200 ;
        RECT 71.000 66.800 71.400 67.200 ;
        RECT 65.400 66.100 65.800 66.500 ;
        RECT 69.400 65.900 69.800 66.300 ;
        RECT 71.800 65.100 72.200 65.500 ;
        RECT 76.600 65.800 77.000 66.200 ;
        RECT 98.200 68.800 98.600 69.200 ;
        RECT 93.400 66.800 93.800 67.200 ;
        RECT 79.800 66.100 80.200 66.500 ;
        RECT 75.000 61.800 75.400 62.200 ;
        RECT 83.800 65.900 84.200 66.300 ;
        RECT 86.200 65.100 86.600 65.500 ;
        RECT 88.600 65.800 89.000 66.200 ;
        RECT 91.800 65.900 92.200 66.300 ;
        RECT 89.400 65.100 89.800 65.500 ;
        RECT 103.000 66.100 103.400 66.500 ;
        RECT 107.000 65.900 107.400 66.300 ;
        RECT 109.400 65.100 109.800 65.500 ;
        RECT 113.400 65.800 113.800 66.200 ;
        RECT 119.000 65.800 119.400 66.200 ;
        RECT 114.200 65.100 114.600 65.500 ;
        RECT 139.800 68.800 140.200 69.200 ;
        RECT 123.000 63.800 123.400 64.200 ;
        RECT 129.400 61.800 129.800 62.200 ;
        RECT 131.000 65.100 131.400 65.500 ;
        RECT 146.200 68.800 146.600 69.200 ;
        RECT 139.800 61.800 140.200 62.200 ;
        RECT 154.200 66.800 154.600 67.200 ;
        RECT 163.800 68.800 164.200 69.200 ;
        RECT 159.800 66.800 160.200 67.200 ;
        RECT 160.600 64.800 161.000 65.200 ;
        RECT 164.600 65.800 165.000 66.200 ;
        RECT 167.000 61.800 167.400 62.200 ;
        RECT 171.800 67.800 172.200 68.200 ;
        RECT 188.600 68.800 189.000 69.200 ;
        RECT 180.600 66.800 181.000 67.200 ;
        RECT 169.400 64.800 169.800 65.200 ;
        RECT 173.400 65.800 173.800 66.200 ;
        RECT 175.800 64.800 176.200 65.200 ;
        RECT 182.200 65.900 182.600 66.300 ;
        RECT 179.800 65.100 180.200 65.500 ;
        RECT 178.200 61.800 178.600 62.200 ;
        RECT 187.000 63.800 187.400 64.200 ;
        RECT 15.800 58.800 16.200 59.200 ;
        RECT 12.600 56.800 13.000 57.200 ;
        RECT 10.200 54.800 10.600 55.200 ;
        RECT 11.000 54.800 11.400 55.200 ;
        RECT 7.800 52.800 8.200 53.200 ;
        RECT 15.000 53.800 15.400 54.200 ;
        RECT 9.400 52.800 9.800 53.200 ;
        RECT 6.200 51.800 6.600 52.200 ;
        RECT 18.200 58.800 18.600 59.200 ;
        RECT 19.800 54.800 20.200 55.200 ;
        RECT 28.600 58.800 29.000 59.200 ;
        RECT 23.000 54.800 23.400 55.200 ;
        RECT 23.800 54.800 24.200 55.200 ;
        RECT 27.800 54.800 28.200 55.200 ;
        RECT 20.600 52.800 21.000 53.200 ;
        RECT 21.400 51.800 21.800 52.200 ;
        RECT 27.800 53.800 28.200 54.200 ;
        RECT 31.100 55.900 31.500 56.300 ;
        RECT 31.700 54.900 32.100 55.300 ;
        RECT 31.100 53.100 31.500 53.500 ;
        RECT 35.000 53.800 35.400 54.200 ;
        RECT 32.600 51.800 33.000 52.200 ;
        RECT 35.800 52.800 36.200 53.200 ;
        RECT 42.200 53.800 42.600 54.200 ;
        RECT 51.800 56.800 52.200 57.200 ;
        RECT 49.400 53.800 49.800 54.200 ;
        RECT 43.000 52.800 43.400 53.200 ;
        RECT 59.000 56.200 59.400 56.600 ;
        RECT 60.600 55.500 61.000 55.900 ;
        RECT 61.400 56.800 61.800 57.200 ;
        RECT 68.600 56.200 69.000 56.600 ;
        RECT 70.200 55.500 70.600 55.900 ;
        RECT 75.800 54.800 76.200 55.200 ;
        RECT 76.600 54.800 77.000 55.200 ;
        RECT 60.600 53.100 61.000 53.500 ;
        RECT 70.200 53.100 70.600 53.500 ;
        RECT 71.000 52.800 71.400 53.200 ;
        RECT 73.400 52.800 73.800 53.200 ;
        RECT 74.200 51.800 74.600 52.200 ;
        RECT 87.800 52.800 88.200 53.200 ;
        RECT 85.400 51.800 85.800 52.200 ;
        RECT 90.200 53.800 90.600 54.200 ;
        RECT 92.600 52.800 93.000 53.200 ;
        RECT 111.000 58.800 111.400 59.200 ;
        RECT 101.400 51.800 101.800 52.200 ;
        RECT 107.800 52.800 108.200 53.200 ;
        RECT 117.400 53.800 117.800 54.200 ;
        RECT 122.200 54.800 122.600 55.200 ;
        RECT 121.400 53.800 121.800 54.200 ;
        RECT 118.200 52.800 118.600 53.200 ;
        RECT 131.800 56.200 132.200 56.600 ;
        RECT 133.400 55.500 133.800 55.900 ;
        RECT 133.400 53.100 133.800 53.500 ;
        RECT 124.600 51.800 125.000 52.200 ;
        RECT 135.000 51.800 135.400 52.200 ;
        RECT 140.600 52.800 141.000 53.200 ;
        RECT 147.000 58.800 147.400 59.200 ;
        RECT 155.000 55.900 155.400 56.300 ;
        RECT 162.200 58.800 162.600 59.200 ;
        RECT 163.000 56.800 163.400 57.200 ;
        RECT 147.800 52.800 148.200 53.200 ;
        RECT 151.800 53.800 152.200 54.200 ;
        RECT 152.600 53.800 153.000 54.200 ;
        RECT 155.000 53.100 155.400 53.500 ;
        RECT 163.800 54.800 164.200 55.200 ;
        RECT 157.400 53.200 157.800 53.600 ;
        RECT 165.400 53.800 165.800 54.200 ;
        RECT 171.800 56.800 172.200 57.200 ;
        RECT 170.200 55.800 170.600 56.200 ;
        RECT 168.600 51.800 169.000 52.200 ;
        RECT 173.400 52.800 173.800 53.200 ;
        RECT 176.600 54.800 177.000 55.200 ;
        RECT 192.600 58.800 193.000 59.200 ;
        RECT 182.200 54.800 182.600 55.200 ;
        RECT 177.400 53.800 177.800 54.200 ;
        RECT 178.200 52.800 178.600 53.200 ;
        RECT 183.000 53.800 183.400 54.200 ;
        RECT 183.800 53.100 184.200 53.500 ;
        RECT 180.600 51.800 181.000 52.200 ;
        RECT 193.400 58.800 193.800 59.200 ;
        RECT 194.200 52.800 194.600 53.200 ;
        RECT 3.000 48.800 3.400 49.200 ;
        RECT 8.600 46.800 9.000 47.200 ;
        RECT 23.800 48.800 24.200 49.200 ;
        RECT 15.800 46.800 16.200 47.200 ;
        RECT 33.400 48.800 33.800 49.200 ;
        RECT 20.600 46.800 21.000 47.200 ;
        RECT 5.400 46.100 5.800 46.500 ;
        RECT 9.400 45.900 9.800 46.300 ;
        RECT 12.600 45.800 13.000 46.200 ;
        RECT 11.800 45.100 12.200 45.500 ;
        RECT 14.200 45.800 14.600 46.200 ;
        RECT 15.000 45.100 15.400 45.500 ;
        RECT 24.600 45.100 25.000 45.500 ;
        RECT 38.200 48.800 38.600 49.200 ;
        RECT 39.000 47.800 39.400 48.200 ;
        RECT 38.200 46.800 38.600 47.200 ;
        RECT 43.800 47.400 44.200 47.800 ;
        RECT 47.800 48.800 48.200 49.200 ;
        RECT 45.400 46.800 45.800 47.200 ;
        RECT 42.200 45.800 42.600 46.200 ;
        RECT 58.200 47.800 58.600 48.200 ;
        RECT 55.800 46.800 56.200 47.200 ;
        RECT 50.200 46.100 50.600 46.500 ;
        RECT 54.200 45.900 54.600 46.300 ;
        RECT 56.600 45.100 57.000 45.500 ;
        RECT 47.800 41.800 48.200 42.200 ;
        RECT 68.600 48.800 69.000 49.200 ;
        RECT 73.400 46.800 73.800 47.200 ;
        RECT 78.200 48.800 78.600 49.200 ;
        RECT 71.000 46.100 71.400 46.500 ;
        RECT 77.400 45.100 77.800 45.500 ;
        RECT 86.200 48.800 86.600 49.200 ;
        RECT 83.000 44.800 83.400 45.200 ;
        RECT 84.600 44.800 85.000 45.200 ;
        RECT 93.400 48.800 93.800 49.200 ;
        RECT 87.800 46.800 88.200 47.200 ;
        RECT 91.800 44.800 92.200 45.200 ;
        RECT 99.800 48.800 100.200 49.200 ;
        RECT 99.000 45.800 99.400 46.200 ;
        RECT 111.800 48.800 112.200 49.200 ;
        RECT 115.000 48.800 115.400 49.200 ;
        RECT 118.200 48.800 118.600 49.200 ;
        RECT 119.800 48.800 120.200 49.200 ;
        RECT 113.400 46.800 113.800 47.200 ;
        RECT 115.800 45.800 116.200 46.200 ;
        RECT 139.000 48.800 139.400 49.200 ;
        RECT 127.800 46.800 128.200 47.200 ;
        RECT 122.200 46.100 122.600 46.500 ;
        RECT 126.200 45.900 126.600 46.300 ;
        RECT 128.600 45.100 129.000 45.500 ;
        RECT 129.400 45.100 129.800 45.500 ;
        RECT 144.600 46.800 145.000 47.200 ;
        RECT 141.400 46.100 141.800 46.500 ;
        RECT 145.400 45.900 145.800 46.300 ;
        RECT 147.800 45.100 148.200 45.500 ;
        RECT 156.600 48.800 157.000 49.200 ;
        RECT 158.200 48.800 158.600 49.200 ;
        RECT 151.800 45.800 152.200 46.200 ;
        RECT 154.200 45.800 154.600 46.200 ;
        RECT 156.600 45.800 157.000 46.200 ;
        RECT 168.600 47.800 169.000 48.200 ;
        RECT 166.200 46.800 166.600 47.200 ;
        RECT 160.600 46.100 161.000 46.500 ;
        RECT 164.600 45.900 165.000 46.300 ;
        RECT 167.000 45.100 167.400 45.500 ;
        RECT 167.800 44.800 168.200 45.200 ;
        RECT 181.400 48.800 181.800 49.200 ;
        RECT 173.400 46.800 173.800 47.200 ;
        RECT 191.000 48.800 191.400 49.200 ;
        RECT 171.800 45.800 172.200 46.200 ;
        RECT 175.000 45.900 175.400 46.300 ;
        RECT 172.600 45.100 173.000 45.500 ;
        RECT 182.200 45.100 182.600 45.500 ;
        RECT 0.600 38.800 1.000 39.200 ;
        RECT 7.800 36.200 8.200 36.600 ;
        RECT 9.400 35.500 9.800 35.900 ;
        RECT 10.200 38.800 10.600 39.200 ;
        RECT 17.400 36.200 17.800 36.600 ;
        RECT 19.000 35.500 19.400 35.900 ;
        RECT 28.600 38.800 29.000 39.200 ;
        RECT 9.400 33.100 9.800 33.500 ;
        RECT 19.000 33.100 19.400 33.500 ;
        RECT 19.800 33.100 20.200 33.500 ;
        RECT 36.600 36.200 37.000 36.600 ;
        RECT 38.200 35.500 38.600 35.900 ;
        RECT 35.800 32.800 36.200 33.200 ;
        RECT 29.400 31.800 29.800 32.200 ;
        RECT 38.200 33.100 38.600 33.500 ;
        RECT 43.000 34.800 43.400 35.200 ;
        RECT 53.400 38.800 53.800 39.200 ;
        RECT 44.600 34.800 45.000 35.200 ;
        RECT 52.600 34.800 53.000 35.200 ;
        RECT 60.600 36.200 61.000 36.600 ;
        RECT 62.200 35.500 62.600 35.900 ;
        RECT 57.400 34.800 57.800 35.200 ;
        RECT 54.200 33.800 54.600 34.200 ;
        RECT 52.600 32.800 53.000 33.200 ;
        RECT 62.200 33.100 62.600 33.500 ;
        RECT 66.200 32.800 66.600 33.200 ;
        RECT 71.800 33.800 72.200 34.200 ;
        RECT 88.600 38.800 89.000 39.200 ;
        RECT 78.200 32.800 78.600 33.200 ;
        RECT 84.600 34.800 85.000 35.200 ;
        RECT 99.800 38.800 100.200 39.200 ;
        RECT 79.800 33.100 80.200 33.500 ;
        RECT 89.400 33.100 89.800 33.500 ;
        RECT 91.800 32.800 92.200 33.200 ;
        RECT 112.600 36.800 113.000 37.200 ;
        RECT 102.200 34.000 102.600 34.400 ;
        RECT 114.200 35.800 114.600 36.200 ;
        RECT 119.800 36.200 120.200 36.600 ;
        RECT 124.600 38.800 125.000 39.200 ;
        RECT 121.400 35.500 121.800 35.900 ;
        RECT 111.800 32.800 112.200 33.200 ;
        RECT 121.400 33.100 121.800 33.500 ;
        RECT 122.200 32.800 122.600 33.200 ;
        RECT 131.800 36.200 132.200 36.600 ;
        RECT 133.400 35.500 133.800 35.900 ;
        RECT 133.400 33.100 133.800 33.500 ;
        RECT 144.600 38.800 145.000 39.200 ;
        RECT 156.600 38.800 157.000 39.200 ;
        RECT 151.000 34.800 151.400 35.200 ;
        RECT 166.200 38.800 166.600 39.200 ;
        RECT 144.600 31.800 145.000 32.200 ;
        RECT 147.800 33.100 148.200 33.500 ;
        RECT 162.200 34.800 162.600 35.200 ;
        RECT 158.200 33.800 158.600 34.200 ;
        RECT 150.200 32.800 150.600 33.200 ;
        RECT 157.400 33.100 157.800 33.500 ;
        RECT 177.400 36.200 177.800 36.600 ;
        RECT 179.000 35.500 179.400 35.900 ;
        RECT 187.000 36.800 187.400 37.200 ;
        RECT 179.000 33.100 179.400 33.500 ;
        RECT 170.200 31.800 170.600 32.200 ;
        RECT 179.800 33.100 180.200 33.500 ;
        RECT 188.600 31.800 189.000 32.200 ;
        RECT 9.400 26.800 9.800 27.200 ;
        RECT 8.600 25.100 9.000 25.500 ;
        RECT 36.600 28.800 37.000 29.200 ;
        RECT 20.600 25.900 21.000 26.300 ;
        RECT 17.400 21.800 17.800 22.200 ;
        RECT 18.200 25.100 18.600 25.500 ;
        RECT 28.600 26.800 29.000 27.200 ;
        RECT 30.200 25.900 30.600 26.300 ;
        RECT 27.000 21.800 27.400 22.200 ;
        RECT 27.800 25.100 28.200 25.500 ;
        RECT 48.600 28.800 49.000 29.200 ;
        RECT 40.600 26.800 41.000 27.200 ;
        RECT 54.200 28.800 54.600 29.200 ;
        RECT 37.400 25.800 37.800 26.200 ;
        RECT 42.200 25.900 42.600 26.300 ;
        RECT 39.800 25.100 40.200 25.500 ;
        RECT 51.000 26.800 51.400 27.200 ;
        RECT 59.800 26.800 60.200 27.200 ;
        RECT 56.600 26.100 57.000 26.500 ;
        RECT 60.600 25.900 61.000 26.300 ;
        RECT 63.000 25.100 63.400 25.500 ;
        RECT 71.800 25.800 72.200 26.200 ;
        RECT 83.800 26.800 84.200 27.200 ;
        RECT 80.600 26.100 81.000 26.500 ;
        RECT 84.600 25.900 85.000 26.300 ;
        RECT 91.800 26.800 92.200 27.200 ;
        RECT 95.800 26.800 96.200 27.200 ;
        RECT 99.000 26.800 99.400 27.200 ;
        RECT 90.200 26.100 90.600 26.500 ;
        RECT 87.000 25.100 87.400 25.500 ;
        RECT 78.200 21.800 78.600 22.200 ;
        RECT 96.600 25.100 97.000 25.500 ;
        RECT 87.800 21.800 88.200 22.200 ;
        RECT 122.200 28.800 122.600 29.200 ;
        RECT 104.600 26.100 105.000 26.500 ;
        RECT 108.600 25.900 109.000 26.300 ;
        RECT 114.200 26.100 114.600 26.500 ;
        RECT 111.000 25.100 111.400 25.500 ;
        RECT 102.200 21.800 102.600 22.200 ;
        RECT 120.600 25.100 121.000 25.500 ;
        RECT 111.800 21.800 112.200 22.200 ;
        RECT 123.800 28.800 124.200 29.200 ;
        RECT 123.800 21.800 124.200 22.200 ;
        RECT 135.000 26.800 135.400 27.200 ;
        RECT 154.200 28.800 154.600 29.200 ;
        RECT 133.400 25.800 133.800 26.200 ;
        RECT 134.200 25.100 134.600 25.500 ;
        RECT 141.400 23.800 141.800 24.200 ;
        RECT 143.000 21.800 143.400 22.200 ;
        RECT 145.400 25.100 145.800 25.500 ;
        RECT 164.600 28.800 165.000 29.200 ;
        RECT 167.800 28.800 168.200 29.200 ;
        RECT 157.400 25.900 157.800 26.300 ;
        RECT 155.000 25.100 155.400 25.500 ;
        RECT 188.600 28.800 189.000 29.200 ;
        RECT 180.600 26.800 181.000 27.200 ;
        RECT 170.200 26.100 170.600 26.500 ;
        RECT 174.200 25.900 174.600 26.300 ;
        RECT 176.600 25.100 177.000 25.500 ;
        RECT 179.000 25.800 179.400 26.200 ;
        RECT 182.200 25.900 182.600 26.300 ;
        RECT 179.800 25.100 180.200 25.500 ;
        RECT 188.600 21.800 189.000 22.200 ;
        RECT 10.200 16.200 10.600 16.600 ;
        RECT 11.800 15.500 12.200 15.900 ;
        RECT 25.400 18.800 25.800 19.200 ;
        RECT 11.800 13.100 12.200 13.500 ;
        RECT 3.000 11.800 3.400 12.200 ;
        RECT 14.200 12.800 14.600 13.200 ;
        RECT 15.000 13.100 15.400 13.500 ;
        RECT 13.400 11.800 13.800 12.200 ;
        RECT 23.800 11.800 24.200 12.200 ;
        RECT 30.200 13.800 30.600 14.200 ;
        RECT 35.000 16.800 35.400 17.200 ;
        RECT 26.200 12.800 26.600 13.200 ;
        RECT 28.600 12.800 29.000 13.200 ;
        RECT 42.200 16.200 42.600 16.600 ;
        RECT 43.800 15.500 44.200 15.900 ;
        RECT 34.200 12.800 34.600 13.200 ;
        RECT 43.800 13.100 44.200 13.500 ;
        RECT 49.400 16.800 49.800 17.200 ;
        RECT 56.600 16.200 57.000 16.600 ;
        RECT 58.200 15.500 58.600 15.900 ;
        RECT 59.800 18.800 60.200 19.200 ;
        RECT 69.400 14.800 69.800 15.200 ;
        RECT 48.600 11.800 49.000 12.200 ;
        RECT 67.000 13.800 67.400 14.200 ;
        RECT 58.200 13.100 58.600 13.500 ;
        RECT 66.200 13.100 66.600 13.500 ;
        RECT 75.800 16.800 76.200 17.200 ;
        RECT 79.000 13.800 79.400 14.200 ;
        RECT 87.800 18.800 88.200 19.200 ;
        RECT 80.600 13.800 81.000 14.200 ;
        RECT 75.000 11.800 75.400 12.200 ;
        RECT 79.800 12.800 80.200 13.200 ;
        RECT 83.000 12.800 83.400 13.200 ;
        RECT 83.800 12.800 84.200 13.200 ;
        RECT 90.200 14.800 90.600 15.200 ;
        RECT 91.000 13.800 91.400 14.200 ;
        RECT 93.400 12.800 93.800 13.200 ;
        RECT 100.600 12.800 101.000 13.200 ;
        RECT 115.800 11.800 116.200 12.200 ;
        RECT 128.600 16.200 129.000 16.600 ;
        RECT 130.200 15.500 130.600 15.900 ;
        RECT 135.000 14.800 135.400 15.200 ;
        RECT 137.400 14.800 137.800 15.200 ;
        RECT 152.600 18.800 153.000 19.200 ;
        RECT 150.200 16.800 150.600 17.200 ;
        RECT 130.200 13.100 130.600 13.500 ;
        RECT 131.000 12.800 131.400 13.200 ;
        RECT 135.800 13.800 136.200 14.200 ;
        RECT 131.800 11.800 132.200 12.200 ;
        RECT 143.000 13.100 143.400 13.500 ;
        RECT 154.200 13.800 154.600 14.200 ;
        RECT 141.400 11.800 141.800 12.200 ;
        RECT 145.400 12.800 145.800 13.200 ;
        RECT 155.000 12.800 155.400 13.200 ;
        RECT 163.000 14.800 163.400 15.200 ;
        RECT 157.400 13.800 157.800 14.200 ;
        RECT 158.200 12.800 158.600 13.200 ;
        RECT 159.000 13.100 159.400 13.500 ;
        RECT 174.200 18.800 174.600 19.200 ;
        RECT 167.800 11.800 168.200 12.200 ;
        RECT 184.600 18.800 185.000 19.200 ;
        RECT 179.800 14.800 180.200 15.200 ;
        RECT 183.000 14.800 183.400 15.200 ;
        RECT 177.400 13.800 177.800 14.200 ;
        RECT 180.600 13.800 181.000 14.200 ;
        RECT 183.000 12.800 183.400 13.200 ;
        RECT 183.800 12.800 184.200 13.200 ;
        RECT 186.200 13.800 186.600 14.200 ;
        RECT 185.400 13.100 185.800 13.500 ;
        RECT 194.200 11.800 194.600 12.200 ;
        RECT 11.800 8.800 12.200 9.200 ;
        RECT 8.600 6.800 9.000 7.200 ;
        RECT 4.600 4.800 5.000 5.200 ;
        RECT 12.600 7.800 13.000 8.200 ;
        RECT 19.000 8.800 19.400 9.200 ;
        RECT 17.400 7.800 17.800 8.200 ;
        RECT 30.200 8.800 30.600 9.200 ;
        RECT 33.400 8.800 33.800 9.200 ;
        RECT 35.000 8.800 35.400 9.200 ;
        RECT 11.800 6.800 12.200 7.200 ;
        RECT 14.200 5.800 14.600 6.200 ;
        RECT 27.000 7.800 27.400 8.200 ;
        RECT 16.600 4.800 17.000 5.200 ;
        RECT 25.400 5.800 25.800 6.200 ;
        RECT 31.000 6.800 31.400 7.200 ;
        RECT 29.400 5.800 29.800 6.200 ;
        RECT 32.600 4.800 33.000 5.200 ;
        RECT 37.400 6.100 37.800 6.500 ;
        RECT 41.400 5.900 41.800 6.300 ;
        RECT 49.400 5.800 49.800 6.200 ;
        RECT 43.800 5.100 44.200 5.500 ;
        RECT 48.600 4.800 49.000 5.200 ;
        RECT 63.800 8.800 64.200 9.200 ;
        RECT 51.000 5.800 51.400 6.200 ;
        RECT 59.800 6.800 60.200 7.200 ;
        RECT 55.800 4.800 56.200 5.200 ;
        RECT 74.200 7.800 74.600 8.200 ;
        RECT 75.000 7.800 75.400 8.200 ;
        RECT 69.400 5.800 69.800 6.200 ;
        RECT 63.800 4.800 64.200 5.200 ;
        RECT 64.600 5.100 65.000 5.500 ;
        RECT 77.400 8.800 77.800 9.200 ;
        RECT 76.600 6.800 77.000 7.200 ;
        RECT 81.400 8.800 81.800 9.200 ;
        RECT 85.400 5.800 85.800 6.200 ;
        RECT 87.000 4.800 87.400 5.200 ;
        RECT 84.600 2.800 85.000 3.200 ;
        RECT 89.400 5.100 89.800 5.500 ;
        RECT 102.200 5.800 102.600 6.200 ;
        RECT 98.200 3.800 98.600 4.200 ;
        RECT 103.000 4.800 103.400 5.200 ;
        RECT 113.400 6.800 113.800 7.200 ;
        RECT 111.000 6.100 111.400 6.500 ;
        RECT 115.000 5.900 115.400 6.300 ;
        RECT 117.400 5.100 117.800 5.500 ;
        RECT 108.600 3.800 109.000 4.200 ;
        RECT 137.400 8.800 137.800 9.200 ;
        RECT 124.600 6.800 125.000 7.200 ;
        RECT 120.600 5.800 121.000 6.200 ;
        RECT 129.400 6.800 129.800 7.200 ;
        RECT 140.600 8.800 141.000 9.200 ;
        RECT 125.400 4.800 125.800 5.200 ;
        RECT 127.800 4.800 128.200 5.200 ;
        RECT 128.600 5.100 129.000 5.500 ;
        RECT 150.200 8.800 150.600 9.200 ;
        RECT 141.400 5.100 141.800 5.500 ;
        RECT 155.000 6.100 155.400 6.500 ;
        RECT 161.400 5.100 161.800 5.500 ;
        RECT 163.800 5.800 164.200 6.200 ;
        RECT 172.600 8.800 173.000 9.200 ;
        RECT 163.000 4.800 163.400 5.200 ;
        RECT 169.400 4.800 169.800 5.200 ;
        RECT 171.800 5.800 172.200 6.200 ;
        RECT 194.200 8.800 194.600 9.200 ;
        RECT 185.400 6.800 185.800 7.200 ;
        RECT 175.000 6.100 175.400 6.500 ;
        RECT 182.200 5.800 182.600 6.200 ;
        RECT 181.400 5.100 181.800 5.500 ;
        RECT 184.600 5.100 185.000 5.500 ;
      LAYER metal2 ;
        RECT 6.200 167.800 6.600 168.200 ;
        RECT 7.000 167.800 7.400 168.200 ;
        RECT 9.400 167.800 9.800 168.200 ;
        RECT 12.600 167.800 13.000 168.200 ;
        RECT 13.400 167.800 13.800 168.200 ;
        RECT 19.800 168.100 20.200 168.200 ;
        RECT 20.600 168.100 21.000 168.200 ;
        RECT 19.800 167.800 21.000 168.100 ;
        RECT 21.400 167.800 21.800 168.200 ;
        RECT 6.200 167.200 6.500 167.800 ;
        RECT 2.200 166.800 2.600 167.200 ;
        RECT 5.400 166.800 5.800 167.200 ;
        RECT 6.200 166.800 6.600 167.200 ;
        RECT 2.200 166.200 2.500 166.800 ;
        RECT 5.400 166.200 5.700 166.800 ;
        RECT 2.200 165.800 2.600 166.200 ;
        RECT 5.400 165.800 5.800 166.200 ;
        RECT 7.000 164.200 7.300 167.800 ;
        RECT 9.400 167.200 9.700 167.800 ;
        RECT 9.400 166.800 9.800 167.200 ;
        RECT 11.000 167.100 11.400 167.200 ;
        RECT 11.800 167.100 12.200 167.200 ;
        RECT 11.000 166.800 12.200 167.100 ;
        RECT 7.800 166.100 8.200 166.200 ;
        RECT 8.600 166.100 9.000 166.200 ;
        RECT 7.800 165.800 9.000 166.100 ;
        RECT 10.200 165.800 10.600 166.200 ;
        RECT 11.800 165.800 12.200 166.200 ;
        RECT 10.200 164.200 10.500 165.800 ;
        RECT 11.800 165.200 12.100 165.800 ;
        RECT 11.800 164.800 12.200 165.200 ;
        RECT 7.000 163.800 7.400 164.200 ;
        RECT 10.200 163.800 10.600 164.200 ;
        RECT 12.600 159.200 12.900 167.800 ;
        RECT 13.400 167.200 13.700 167.800 ;
        RECT 13.400 166.800 13.800 167.200 ;
        RECT 14.200 166.800 14.600 167.200 ;
        RECT 18.200 166.800 18.600 167.200 ;
        RECT 14.200 164.200 14.500 166.800 ;
        RECT 18.200 166.200 18.500 166.800 ;
        RECT 15.000 165.800 15.400 166.200 ;
        RECT 15.800 166.100 16.200 166.200 ;
        RECT 16.600 166.100 17.000 166.200 ;
        RECT 15.800 165.800 17.000 166.100 ;
        RECT 18.200 165.800 18.600 166.200 ;
        RECT 15.000 165.200 15.300 165.800 ;
        RECT 15.000 164.800 15.400 165.200 ;
        RECT 14.200 163.800 14.600 164.200 ;
        RECT 12.600 158.800 13.000 159.200 ;
        RECT 0.600 151.800 1.000 152.200 ;
        RECT 3.000 152.100 3.400 157.900 ;
        RECT 6.200 154.800 6.600 155.200 ;
        RECT 0.600 144.200 0.900 151.800 ;
        RECT 0.600 144.100 1.000 144.200 ;
        RECT 1.400 144.100 1.800 144.200 ;
        RECT 0.600 143.800 1.800 144.100 ;
        RECT 3.000 143.100 3.400 148.900 ;
        RECT 6.200 147.200 6.500 154.800 ;
        RECT 7.000 152.800 7.400 153.200 ;
        RECT 6.200 146.800 6.600 147.200 ;
        RECT 6.200 146.200 6.500 146.800 ;
        RECT 6.200 145.800 6.600 146.200 ;
        RECT 7.000 140.200 7.300 152.800 ;
        RECT 7.800 152.100 8.200 157.900 ;
        RECT 9.400 153.100 9.800 155.900 ;
        RECT 10.200 154.800 10.600 155.200 ;
        RECT 14.200 154.800 14.600 155.200 ;
        RECT 7.800 143.100 8.200 148.900 ;
        RECT 8.600 146.800 9.000 147.200 ;
        RECT 7.000 139.800 7.400 140.200 ;
        RECT 0.600 136.800 1.000 137.200 ;
        RECT 0.600 136.200 0.900 136.800 ;
        RECT 0.600 135.800 1.000 136.200 ;
        RECT 3.000 132.100 3.400 137.900 ;
        RECT 6.200 134.800 6.600 135.200 ;
        RECT 6.200 134.200 6.500 134.800 ;
        RECT 7.000 134.200 7.300 139.800 ;
        RECT 6.200 133.800 6.600 134.200 ;
        RECT 7.000 133.800 7.400 134.200 ;
        RECT 6.200 129.800 6.600 130.200 ;
        RECT 0.600 124.100 1.000 124.200 ;
        RECT 1.400 124.100 1.800 124.200 ;
        RECT 0.600 123.800 1.800 124.100 ;
        RECT 0.600 119.200 0.900 123.800 ;
        RECT 3.000 123.100 3.400 128.900 ;
        RECT 6.200 126.200 6.500 129.800 ;
        RECT 6.200 125.800 6.600 126.200 ;
        RECT 0.600 118.800 1.000 119.200 ;
        RECT 3.000 112.100 3.400 117.900 ;
        RECT 6.200 115.200 6.500 125.800 ;
        RECT 6.200 114.800 6.600 115.200 ;
        RECT 7.000 114.200 7.300 133.800 ;
        RECT 7.800 132.100 8.200 137.900 ;
        RECT 7.800 123.100 8.200 128.900 ;
        RECT 8.600 128.200 8.900 146.800 ;
        RECT 9.400 145.100 9.800 147.900 ;
        RECT 10.200 145.100 10.500 154.800 ;
        RECT 14.200 154.200 14.500 154.800 ;
        RECT 15.000 154.200 15.300 164.800 ;
        RECT 21.400 159.200 21.700 167.800 ;
        RECT 25.400 163.100 25.800 168.900 ;
        RECT 29.400 165.900 29.800 166.300 ;
        RECT 29.400 165.200 29.700 165.900 ;
        RECT 29.400 164.800 29.800 165.200 ;
        RECT 26.200 163.800 26.600 164.200 ;
        RECT 23.000 162.100 23.400 162.200 ;
        RECT 23.800 162.100 24.200 162.200 ;
        RECT 23.000 161.800 24.200 162.100 ;
        RECT 25.400 161.800 25.800 162.200 ;
        RECT 21.400 158.800 21.800 159.200 ;
        RECT 25.400 155.200 25.700 161.800 ;
        RECT 26.200 159.200 26.500 163.800 ;
        RECT 30.200 163.100 30.600 168.900 ;
        RECT 31.000 166.800 31.400 167.200 ;
        RECT 26.200 158.800 26.600 159.200 ;
        RECT 31.000 157.200 31.300 166.800 ;
        RECT 31.800 165.100 32.200 167.900 ;
        RECT 35.000 163.100 35.400 168.900 ;
        RECT 39.000 165.900 39.400 166.300 ;
        RECT 39.000 165.200 39.300 165.900 ;
        RECT 39.000 164.800 39.400 165.200 ;
        RECT 39.800 163.100 40.200 168.900 ;
        RECT 40.600 167.800 41.000 168.200 ;
        RECT 42.200 168.100 42.600 168.200 ;
        RECT 43.000 168.100 43.400 168.200 ;
        RECT 40.600 167.200 40.900 167.800 ;
        RECT 40.600 166.800 41.000 167.200 ;
        RECT 41.400 165.100 41.800 167.900 ;
        RECT 42.200 167.800 43.400 168.100 ;
        RECT 31.800 162.100 32.200 162.200 ;
        RECT 32.600 162.100 33.000 162.200 ;
        RECT 31.800 161.800 33.000 162.100 ;
        RECT 31.000 156.800 31.400 157.200 ;
        RECT 15.800 154.800 16.200 155.200 ;
        RECT 16.600 154.800 17.000 155.200 ;
        RECT 19.000 154.800 19.400 155.200 ;
        RECT 19.800 155.100 20.200 155.200 ;
        RECT 20.600 155.100 21.000 155.200 ;
        RECT 19.800 154.800 21.000 155.100 ;
        RECT 23.800 154.800 24.200 155.200 ;
        RECT 25.400 154.800 25.800 155.200 ;
        RECT 28.600 154.800 29.000 155.200 ;
        RECT 14.200 153.800 14.600 154.200 ;
        RECT 15.000 153.800 15.400 154.200 ;
        RECT 11.000 146.800 11.400 147.200 ;
        RECT 11.800 146.800 12.200 147.200 ;
        RECT 11.000 146.200 11.300 146.800 ;
        RECT 11.800 146.200 12.100 146.800 ;
        RECT 11.000 145.800 11.400 146.200 ;
        RECT 11.800 145.800 12.200 146.200 ;
        RECT 12.600 145.800 13.000 146.200 ;
        RECT 13.400 145.800 13.800 146.200 ;
        RECT 14.200 146.100 14.600 146.200 ;
        RECT 15.000 146.100 15.400 146.200 ;
        RECT 14.200 145.800 15.400 146.100 ;
        RECT 10.200 144.800 11.300 145.100 ;
        RECT 9.400 133.100 9.800 135.900 ;
        RECT 10.200 133.100 10.600 135.900 ;
        RECT 8.600 127.800 9.000 128.200 ;
        RECT 8.600 127.200 8.900 127.800 ;
        RECT 8.600 126.800 9.000 127.200 ;
        RECT 9.400 125.100 9.800 127.900 ;
        RECT 11.000 127.200 11.300 144.800 ;
        RECT 11.800 132.100 12.200 137.900 ;
        RECT 12.600 135.200 12.900 145.800 ;
        RECT 13.400 144.200 13.700 145.800 ;
        RECT 13.400 143.800 13.800 144.200 ;
        RECT 15.800 137.200 16.100 154.800 ;
        RECT 16.600 146.200 16.900 154.800 ;
        RECT 19.000 154.200 19.300 154.800 ;
        RECT 19.000 153.800 19.400 154.200 ;
        RECT 20.600 151.200 20.900 154.800 ;
        RECT 23.800 154.200 24.100 154.800 ;
        RECT 23.800 153.800 24.200 154.200 ;
        RECT 20.600 150.800 21.000 151.200 ;
        RECT 16.600 145.800 17.000 146.200 ;
        RECT 19.800 143.100 20.200 148.900 ;
        RECT 23.800 147.800 24.200 148.200 ;
        RECT 23.800 146.300 24.100 147.800 ;
        RECT 20.600 145.800 21.000 146.200 ;
        RECT 23.800 145.900 24.200 146.300 ;
        RECT 17.400 142.100 17.800 142.200 ;
        RECT 18.200 142.100 18.600 142.200 ;
        RECT 17.400 141.800 18.600 142.100 ;
        RECT 15.800 136.800 16.200 137.200 ;
        RECT 12.600 134.800 13.000 135.200 ;
        RECT 13.400 134.800 13.800 135.200 ;
        RECT 13.400 134.200 13.700 134.800 ;
        RECT 13.400 133.800 13.800 134.200 ;
        RECT 14.200 133.800 14.600 134.200 ;
        RECT 14.200 133.200 14.500 133.800 ;
        RECT 14.200 132.800 14.600 133.200 ;
        RECT 11.000 126.800 11.400 127.200 ;
        RECT 8.600 123.800 9.000 124.200 ;
        RECT 7.000 113.800 7.400 114.200 ;
        RECT 7.800 112.100 8.200 117.900 ;
        RECT 8.600 108.200 8.900 123.800 ;
        RECT 12.600 123.100 13.000 128.900 ;
        RECT 14.200 127.200 14.500 132.800 ;
        RECT 14.200 126.800 14.600 127.200 ;
        RECT 15.800 126.200 16.100 136.800 ;
        RECT 16.600 132.100 17.000 137.900 ;
        RECT 19.000 136.800 19.400 137.200 ;
        RECT 19.000 136.200 19.300 136.800 ;
        RECT 19.000 135.800 19.400 136.200 ;
        RECT 19.800 134.800 20.200 135.200 ;
        RECT 19.800 134.200 20.100 134.800 ;
        RECT 19.800 133.800 20.200 134.200 ;
        RECT 20.600 133.200 20.900 145.800 ;
        RECT 24.600 143.100 25.000 148.900 ;
        RECT 25.400 146.200 25.700 154.800 ;
        RECT 28.600 154.200 28.900 154.800 ;
        RECT 28.600 153.800 29.000 154.200 ;
        RECT 29.400 152.100 29.800 152.200 ;
        RECT 30.200 152.100 30.600 152.200 ;
        RECT 31.800 152.100 32.200 157.900 ;
        RECT 35.800 155.800 36.200 156.200 ;
        RECT 35.800 155.100 36.100 155.800 ;
        RECT 35.800 154.700 36.200 155.100 ;
        RECT 32.600 153.800 33.000 154.200 ;
        RECT 29.400 151.800 30.600 152.100 ;
        RECT 31.000 149.800 31.400 150.200 ;
        RECT 25.400 145.800 25.800 146.200 ;
        RECT 25.400 142.100 25.700 145.800 ;
        RECT 26.200 145.100 26.600 147.900 ;
        RECT 28.600 143.800 29.000 144.200 ;
        RECT 25.400 141.800 26.500 142.100 ;
        RECT 25.400 139.800 25.800 140.200 ;
        RECT 23.000 135.800 23.400 136.200 ;
        RECT 23.000 135.200 23.300 135.800 ;
        RECT 21.400 134.800 21.800 135.200 ;
        RECT 22.200 134.800 22.600 135.200 ;
        RECT 23.000 134.800 23.400 135.200 ;
        RECT 21.400 133.200 21.700 134.800 ;
        RECT 22.200 134.200 22.500 134.800 ;
        RECT 22.200 133.800 22.600 134.200 ;
        RECT 19.000 133.100 19.400 133.200 ;
        RECT 19.800 133.100 20.200 133.200 ;
        RECT 19.000 132.800 20.200 133.100 ;
        RECT 20.600 132.800 21.000 133.200 ;
        RECT 21.400 132.800 21.800 133.200 ;
        RECT 16.600 126.800 17.000 127.200 ;
        RECT 16.600 126.300 16.900 126.800 ;
        RECT 15.800 125.800 16.200 126.200 ;
        RECT 16.600 125.900 17.000 126.300 ;
        RECT 17.400 123.100 17.800 128.900 ;
        RECT 18.200 126.800 18.600 127.200 ;
        RECT 10.200 121.800 10.600 122.200 ;
        RECT 10.200 117.200 10.500 121.800 ;
        RECT 10.200 116.800 10.600 117.200 ;
        RECT 9.400 113.100 9.800 115.900 ;
        RECT 11.800 115.100 12.200 115.200 ;
        RECT 12.600 115.100 13.000 115.200 ;
        RECT 11.800 114.800 13.000 115.100 ;
        RECT 13.400 114.800 13.800 115.200 ;
        RECT 13.400 114.400 13.700 114.800 ;
        RECT 13.400 114.300 13.800 114.400 ;
        RECT 14.200 114.300 14.600 114.400 ;
        RECT 10.200 113.800 10.600 114.200 ;
        RECT 11.800 114.100 12.200 114.200 ;
        RECT 12.600 114.100 13.000 114.200 ;
        RECT 11.800 113.800 13.000 114.100 ;
        RECT 13.400 114.000 14.600 114.300 ;
        RECT 13.400 113.800 13.700 114.000 ;
        RECT 10.200 113.200 10.500 113.800 ;
        RECT 10.200 112.800 10.600 113.200 ;
        RECT 15.800 113.100 16.200 115.900 ;
        RECT 11.000 111.800 11.400 112.200 ;
        RECT 15.000 111.800 15.400 112.200 ;
        RECT 17.400 112.100 17.800 117.900 ;
        RECT 18.200 113.200 18.500 126.800 ;
        RECT 19.000 125.100 19.400 127.900 ;
        RECT 19.800 125.100 20.200 127.900 ;
        RECT 21.400 123.100 21.800 128.900 ;
        RECT 19.000 114.800 19.400 115.200 ;
        RECT 19.000 113.200 19.300 114.800 ;
        RECT 18.200 112.800 18.600 113.200 ;
        RECT 19.000 112.800 19.400 113.200 ;
        RECT 11.000 109.200 11.300 111.800 ;
        RECT 11.000 108.800 11.400 109.200 ;
        RECT 15.000 108.200 15.300 111.800 ;
        RECT 15.800 108.800 16.200 109.200 ;
        RECT 7.000 108.100 7.400 108.200 ;
        RECT 7.800 108.100 8.200 108.200 ;
        RECT 7.000 107.800 8.200 108.100 ;
        RECT 8.600 107.800 9.000 108.200 ;
        RECT 11.000 107.800 11.400 108.200 ;
        RECT 12.600 107.800 13.000 108.200 ;
        RECT 15.000 107.800 15.400 108.200 ;
        RECT 0.600 107.100 1.000 107.200 ;
        RECT 1.400 107.100 1.800 107.200 ;
        RECT 0.600 106.800 1.800 107.100 ;
        RECT 7.800 106.800 8.200 107.200 ;
        RECT 8.600 107.000 8.900 107.800 ;
        RECT 11.000 107.200 11.300 107.800 ;
        RECT 5.400 105.800 5.800 106.200 ;
        RECT 2.200 104.800 2.600 105.200 ;
        RECT 2.200 104.200 2.500 104.800 ;
        RECT 5.400 104.200 5.700 105.800 ;
        RECT 2.200 103.800 2.600 104.200 ;
        RECT 5.400 103.800 5.800 104.200 ;
        RECT 1.400 95.800 1.800 96.200 ;
        RECT 2.200 96.100 2.600 96.200 ;
        RECT 3.000 96.100 3.400 96.200 ;
        RECT 2.200 95.800 3.400 96.100 ;
        RECT 1.400 89.200 1.700 95.800 ;
        RECT 5.400 95.200 5.700 103.800 ;
        RECT 2.200 95.100 2.600 95.200 ;
        RECT 3.000 95.100 3.400 95.200 ;
        RECT 2.200 94.800 3.400 95.100 ;
        RECT 5.400 94.800 5.800 95.200 ;
        RECT 3.800 90.800 4.200 91.200 ;
        RECT 2.200 89.800 2.600 90.200 ;
        RECT 1.400 88.800 1.800 89.200 ;
        RECT 0.600 87.100 1.000 87.200 ;
        RECT 1.400 87.100 1.800 87.200 ;
        RECT 0.600 86.800 1.800 87.100 ;
        RECT 2.200 85.200 2.500 89.800 ;
        RECT 3.800 86.200 4.100 90.800 ;
        RECT 5.400 90.200 5.700 94.800 ;
        RECT 7.800 94.200 8.100 106.800 ;
        RECT 8.600 106.600 9.000 107.000 ;
        RECT 11.000 106.800 11.400 107.200 ;
        RECT 12.600 106.200 12.900 107.800 ;
        RECT 13.400 106.800 13.800 107.200 ;
        RECT 13.400 106.200 13.700 106.800 ;
        RECT 15.800 106.200 16.100 108.800 ;
        RECT 16.600 107.800 17.000 108.200 ;
        RECT 17.400 107.800 17.800 108.200 ;
        RECT 16.600 107.200 16.900 107.800 ;
        RECT 17.400 107.200 17.700 107.800 ;
        RECT 16.600 106.800 17.000 107.200 ;
        RECT 17.400 106.800 17.800 107.200 ;
        RECT 10.200 106.100 10.600 106.200 ;
        RECT 11.000 106.100 11.400 106.200 ;
        RECT 10.200 105.800 11.400 106.100 ;
        RECT 12.600 105.800 13.000 106.200 ;
        RECT 13.400 105.800 13.800 106.200 ;
        RECT 14.200 105.800 14.600 106.200 ;
        RECT 15.800 105.800 16.200 106.200 ;
        RECT 14.200 105.200 14.500 105.800 ;
        RECT 12.600 104.800 13.000 105.200 ;
        RECT 14.200 104.800 14.600 105.200 ;
        RECT 12.600 104.200 12.900 104.800 ;
        RECT 12.600 103.800 13.000 104.200 ;
        RECT 15.000 102.100 15.400 102.200 ;
        RECT 15.800 102.100 16.200 102.200 ;
        RECT 15.000 101.800 16.200 102.100 ;
        RECT 13.400 99.100 13.800 99.200 ;
        RECT 14.200 99.100 14.600 99.200 ;
        RECT 13.400 98.800 14.600 99.100 ;
        RECT 8.700 95.900 9.100 96.300 ;
        RECT 11.800 95.900 12.200 96.300 ;
        RECT 7.000 94.100 7.400 94.200 ;
        RECT 6.200 93.800 7.400 94.100 ;
        RECT 7.800 93.800 8.200 94.200 ;
        RECT 5.400 89.800 5.800 90.200 ;
        RECT 6.200 87.200 6.500 93.800 ;
        RECT 8.700 93.500 9.000 95.900 ;
        RECT 9.300 94.900 9.700 95.300 ;
        RECT 9.400 94.200 9.700 94.900 ;
        RECT 11.900 94.200 12.200 95.900 ;
        RECT 9.400 93.900 12.200 94.200 ;
        RECT 9.400 93.500 9.800 93.600 ;
        RECT 11.100 93.500 11.500 93.600 ;
        RECT 11.900 93.500 12.200 93.900 ;
        RECT 8.700 93.200 11.500 93.500 ;
        RECT 7.000 93.100 7.400 93.200 ;
        RECT 7.800 93.100 8.200 93.200 ;
        RECT 8.700 93.100 9.100 93.200 ;
        RECT 11.800 93.100 12.200 93.500 ;
        RECT 12.600 93.800 13.000 94.200 ;
        RECT 12.600 93.200 12.900 93.800 ;
        RECT 7.000 92.800 8.200 93.100 ;
        RECT 12.600 92.800 13.000 93.200 ;
        RECT 8.600 91.800 9.000 92.200 ;
        RECT 10.200 92.100 10.600 92.200 ;
        RECT 11.000 92.100 11.400 92.200 ;
        RECT 10.200 91.800 11.400 92.100 ;
        RECT 6.200 86.800 6.600 87.200 ;
        RECT 6.200 86.200 6.500 86.800 ;
        RECT 8.600 86.200 8.900 91.800 ;
        RECT 11.800 90.800 12.200 91.200 ;
        RECT 11.800 86.200 12.100 90.800 ;
        RECT 12.600 89.200 12.900 92.800 ;
        RECT 15.800 92.100 16.200 97.900 ;
        RECT 16.600 94.800 17.000 95.200 ;
        RECT 13.400 89.800 13.800 90.200 ;
        RECT 12.600 88.800 13.000 89.200 ;
        RECT 3.800 85.800 4.200 86.200 ;
        RECT 6.200 85.800 6.600 86.200 ;
        RECT 7.800 85.800 8.200 86.200 ;
        RECT 8.600 85.800 9.000 86.200 ;
        RECT 11.800 85.800 12.200 86.200 ;
        RECT 2.200 84.800 2.600 85.200 ;
        RECT 5.400 81.800 5.800 82.200 ;
        RECT 5.400 75.200 5.700 81.800 ;
        RECT 6.200 79.200 6.500 85.800 ;
        RECT 7.800 85.200 8.100 85.800 ;
        RECT 7.800 84.800 8.200 85.200 ;
        RECT 10.200 81.800 10.600 82.200 ;
        RECT 10.200 80.200 10.500 81.800 ;
        RECT 10.200 79.800 10.600 80.200 ;
        RECT 11.800 79.800 12.200 80.200 ;
        RECT 6.200 78.800 6.600 79.200 ;
        RECT 9.400 79.100 9.800 79.200 ;
        RECT 10.200 79.100 10.600 79.200 ;
        RECT 9.400 78.800 10.600 79.100 ;
        RECT 5.400 74.800 5.800 75.200 ;
        RECT 7.000 75.100 7.400 75.200 ;
        RECT 7.800 75.100 8.200 75.200 ;
        RECT 7.000 74.800 8.200 75.100 ;
        RECT 9.400 74.800 9.800 75.200 ;
        RECT 9.400 74.200 9.700 74.800 ;
        RECT 7.000 74.100 7.400 74.200 ;
        RECT 7.800 74.100 8.200 74.200 ;
        RECT 7.000 73.800 8.200 74.100 ;
        RECT 9.400 73.800 9.800 74.200 ;
        RECT 9.400 72.800 9.800 73.200 ;
        RECT 9.400 67.200 9.700 72.800 ;
        RECT 10.200 71.800 10.600 72.200 ;
        RECT 10.200 69.200 10.500 71.800 ;
        RECT 10.200 68.800 10.600 69.200 ;
        RECT 9.400 66.800 9.800 67.200 ;
        RECT 8.600 61.800 9.000 62.200 ;
        RECT 7.800 53.100 8.200 53.200 ;
        RECT 8.600 53.100 8.900 61.800 ;
        RECT 9.400 56.800 9.800 57.200 ;
        RECT 9.400 55.200 9.700 56.800 ;
        RECT 10.200 55.800 10.600 56.200 ;
        RECT 10.200 55.200 10.500 55.800 ;
        RECT 9.400 54.800 9.800 55.200 ;
        RECT 10.200 54.800 10.600 55.200 ;
        RECT 11.000 54.800 11.400 55.200 ;
        RECT 11.000 54.200 11.300 54.800 ;
        RECT 11.000 53.800 11.400 54.200 ;
        RECT 7.800 52.800 8.900 53.100 ;
        RECT 6.200 51.800 6.600 52.200 ;
        RECT 3.000 49.100 3.400 49.200 ;
        RECT 3.800 49.100 4.200 49.200 ;
        RECT 3.000 48.800 4.200 49.100 ;
        RECT 5.400 43.100 5.800 48.900 ;
        RECT 0.600 39.100 1.000 39.200 ;
        RECT 1.400 39.100 1.800 39.200 ;
        RECT 0.600 38.800 1.800 39.100 ;
        RECT 3.000 32.100 3.400 37.900 ;
        RECT 6.200 30.200 6.500 51.800 ;
        RECT 8.600 48.200 8.900 52.800 ;
        RECT 9.400 52.800 9.800 53.200 ;
        RECT 8.600 47.800 9.000 48.200 ;
        RECT 8.600 47.200 8.900 47.800 ;
        RECT 8.600 46.800 9.000 47.200 ;
        RECT 7.000 35.800 7.400 36.200 ;
        RECT 7.000 35.100 7.300 35.800 ;
        RECT 7.000 34.700 7.400 35.100 ;
        RECT 7.800 32.100 8.200 37.900 ;
        RECT 8.600 34.200 8.900 46.800 ;
        RECT 9.400 46.300 9.700 52.800 ;
        RECT 11.000 49.200 11.300 53.800 ;
        RECT 9.400 45.900 9.800 46.300 ;
        RECT 9.400 40.200 9.700 45.900 ;
        RECT 10.200 43.100 10.600 48.900 ;
        RECT 11.000 48.800 11.400 49.200 ;
        RECT 11.800 49.100 12.100 79.800 ;
        RECT 12.600 72.100 13.000 77.900 ;
        RECT 12.600 63.100 13.000 68.900 ;
        RECT 12.600 56.800 13.000 57.200 ;
        RECT 12.600 56.200 12.900 56.800 ;
        RECT 12.600 55.800 13.000 56.200 ;
        RECT 13.400 55.200 13.700 89.800 ;
        RECT 15.000 83.100 15.400 88.900 ;
        RECT 16.600 82.200 16.900 94.800 ;
        RECT 18.200 94.200 18.500 112.800 ;
        RECT 22.200 112.100 22.600 117.900 ;
        RECT 23.000 107.100 23.300 134.800 ;
        RECT 23.800 133.100 24.200 133.200 ;
        RECT 24.600 133.100 25.000 133.200 ;
        RECT 23.800 132.800 25.000 133.100 ;
        RECT 23.800 131.800 24.200 132.200 ;
        RECT 23.800 126.200 24.100 131.800 ;
        RECT 25.400 126.200 25.700 139.800 ;
        RECT 26.200 135.200 26.500 141.800 ;
        RECT 27.000 141.800 27.400 142.200 ;
        RECT 27.000 136.200 27.300 141.800 ;
        RECT 28.600 140.200 28.900 143.800 ;
        RECT 29.400 143.100 29.800 148.900 ;
        RECT 28.600 139.800 29.000 140.200 ;
        RECT 27.000 135.800 27.400 136.200 ;
        RECT 26.200 134.800 26.600 135.200 ;
        RECT 29.400 135.100 29.800 135.200 ;
        RECT 30.200 135.100 30.600 135.200 ;
        RECT 29.400 134.800 30.600 135.100 ;
        RECT 31.000 133.200 31.300 149.800 ;
        RECT 32.600 147.200 32.900 153.800 ;
        RECT 36.600 152.100 37.000 157.900 ;
        RECT 37.400 155.800 37.800 156.200 ;
        RECT 37.400 154.200 37.700 155.800 ;
        RECT 37.400 153.800 37.800 154.200 ;
        RECT 38.200 153.100 38.600 155.900 ;
        RECT 39.000 153.100 39.400 155.900 ;
        RECT 40.600 152.100 41.000 157.900 ;
        RECT 41.400 154.700 41.800 155.200 ;
        RECT 41.400 151.100 41.700 154.700 ;
        RECT 40.600 150.800 41.700 151.100 ;
        RECT 42.200 154.200 42.500 167.800 ;
        RECT 43.000 166.800 43.400 167.200 ;
        RECT 43.800 166.800 44.200 167.200 ;
        RECT 43.000 166.200 43.300 166.800 ;
        RECT 43.800 166.200 44.100 166.800 ;
        RECT 43.000 165.800 43.400 166.200 ;
        RECT 43.800 165.800 44.200 166.200 ;
        RECT 44.600 165.800 45.000 166.200 ;
        RECT 47.000 165.800 47.400 166.200 ;
        RECT 47.800 166.100 48.200 166.200 ;
        RECT 48.600 166.100 49.000 166.200 ;
        RECT 47.800 165.800 49.000 166.100 ;
        RECT 49.400 165.800 49.800 166.200 ;
        RECT 44.600 158.200 44.900 165.800 ;
        RECT 47.000 162.200 47.300 165.800 ;
        RECT 49.400 165.200 49.700 165.800 ;
        RECT 49.400 164.800 49.800 165.200 ;
        RECT 53.400 163.100 53.800 168.900 ;
        RECT 57.400 166.800 57.800 167.200 ;
        RECT 57.400 166.300 57.700 166.800 ;
        RECT 55.000 165.800 55.400 166.200 ;
        RECT 57.400 165.900 57.800 166.300 ;
        RECT 47.000 161.800 47.400 162.200 ;
        RECT 51.000 162.100 51.400 162.200 ;
        RECT 51.800 162.100 52.200 162.200 ;
        RECT 51.000 161.800 52.200 162.100 ;
        RECT 44.600 157.800 45.000 158.200 ;
        RECT 42.200 153.800 42.600 154.200 ;
        RECT 40.600 149.200 40.900 150.800 ;
        RECT 42.200 150.200 42.500 153.800 ;
        RECT 43.000 151.800 43.400 152.200 ;
        RECT 45.400 152.100 45.800 157.900 ;
        RECT 51.000 153.800 51.400 154.200 ;
        RECT 51.000 153.200 51.300 153.800 ;
        RECT 51.000 152.800 51.400 153.200 ;
        RECT 47.000 152.100 47.400 152.200 ;
        RECT 47.800 152.100 48.200 152.200 ;
        RECT 47.000 151.800 48.200 152.100 ;
        RECT 42.200 149.800 42.600 150.200 ;
        RECT 33.400 147.800 33.800 148.200 ;
        RECT 32.600 146.800 33.000 147.200 ;
        RECT 33.400 146.300 33.700 147.800 ;
        RECT 33.400 145.900 33.800 146.300 ;
        RECT 34.200 143.100 34.600 148.900 ;
        RECT 40.600 148.800 41.000 149.200 ;
        RECT 35.800 145.100 36.200 147.900 ;
        RECT 39.800 147.800 40.200 148.200 ;
        RECT 39.800 147.200 40.100 147.800 ;
        RECT 43.000 147.200 43.300 151.800 ;
        RECT 51.000 150.200 51.300 152.800 ;
        RECT 51.800 152.100 52.200 152.200 ;
        RECT 52.600 152.100 53.000 152.200 ;
        RECT 54.200 152.100 54.600 157.900 ;
        RECT 55.000 156.200 55.300 165.800 ;
        RECT 58.200 163.100 58.600 168.900 ;
        RECT 59.800 165.100 60.200 167.900 ;
        RECT 62.200 167.800 62.600 168.200 ;
        RECT 62.200 167.200 62.500 167.800 ;
        RECT 62.200 166.800 62.600 167.200 ;
        RECT 60.600 165.800 61.000 166.200 ;
        RECT 61.400 166.100 61.800 166.200 ;
        RECT 62.200 166.100 62.600 166.200 ;
        RECT 61.400 165.800 62.600 166.100 ;
        RECT 60.600 164.200 60.900 165.800 ;
        RECT 60.600 163.800 61.000 164.200 ;
        RECT 64.600 163.800 65.000 164.200 ;
        RECT 63.000 161.800 63.400 162.200 ;
        RECT 56.600 158.800 57.000 159.200 ;
        RECT 55.000 155.800 55.400 156.200 ;
        RECT 55.000 155.200 55.300 155.800 ;
        RECT 55.000 154.800 55.400 155.200 ;
        RECT 51.800 151.800 53.000 152.100 ;
        RECT 56.600 151.200 56.900 158.800 ;
        RECT 57.400 154.800 57.800 155.200 ;
        RECT 57.400 151.200 57.700 154.800 ;
        RECT 58.200 151.800 58.600 152.200 ;
        RECT 59.000 152.100 59.400 157.900 ;
        RECT 59.800 153.800 60.200 154.200 ;
        RECT 59.800 153.200 60.100 153.800 ;
        RECT 59.800 152.800 60.200 153.200 ;
        RECT 60.600 153.100 61.000 155.900 ;
        RECT 60.600 152.100 61.000 152.200 ;
        RECT 61.400 152.100 61.800 152.200 ;
        RECT 60.600 151.800 61.800 152.100 ;
        RECT 56.600 150.800 57.000 151.200 ;
        RECT 57.400 150.800 57.800 151.200 ;
        RECT 51.000 149.800 51.400 150.200 ;
        RECT 53.400 148.800 53.800 149.200 ;
        RECT 53.400 148.200 53.700 148.800 ;
        RECT 47.000 147.500 47.400 147.900 ;
        RECT 47.700 147.500 49.800 147.800 ;
        RECT 50.300 147.500 50.700 147.900 ;
        RECT 53.400 147.800 53.800 148.200 ;
        RECT 36.600 147.100 37.000 147.200 ;
        RECT 37.400 147.100 37.800 147.200 ;
        RECT 36.600 146.800 37.800 147.100 ;
        RECT 39.000 146.800 39.400 147.200 ;
        RECT 39.800 146.800 40.200 147.200 ;
        RECT 41.400 146.800 41.800 147.200 ;
        RECT 42.200 147.100 42.600 147.200 ;
        RECT 43.000 147.100 43.400 147.200 ;
        RECT 42.200 146.800 43.400 147.100 ;
        RECT 43.800 146.800 44.200 147.200 ;
        RECT 47.000 147.100 47.300 147.500 ;
        RECT 47.700 147.400 48.100 147.500 ;
        RECT 49.400 147.400 49.800 147.500 ;
        RECT 47.000 146.800 49.400 147.100 ;
        RECT 37.400 146.100 37.800 146.200 ;
        RECT 38.200 146.100 38.600 146.200 ;
        RECT 37.400 145.800 38.600 146.100 ;
        RECT 36.600 145.100 37.000 145.200 ;
        RECT 37.400 145.100 37.800 145.200 ;
        RECT 36.600 144.800 37.800 145.100 ;
        RECT 35.800 138.800 36.200 139.200 ;
        RECT 35.800 135.200 36.100 138.800 ;
        RECT 36.600 136.200 36.900 144.800 ;
        RECT 39.000 144.200 39.300 146.800 ;
        RECT 41.400 146.200 41.700 146.800 ;
        RECT 41.400 145.800 41.800 146.200 ;
        RECT 42.200 145.800 42.600 146.200 ;
        RECT 42.200 144.200 42.500 145.800 ;
        RECT 39.000 143.800 39.400 144.200 ;
        RECT 42.200 143.800 42.600 144.200 ;
        RECT 38.200 142.800 38.600 143.200 ;
        RECT 38.200 137.200 38.500 142.800 ;
        RECT 38.200 136.800 38.600 137.200 ;
        RECT 36.600 135.800 37.000 136.200 ;
        RECT 31.800 134.800 32.200 135.200 ;
        RECT 32.600 134.800 33.000 135.200 ;
        RECT 35.000 135.100 35.400 135.200 ;
        RECT 34.200 134.800 35.400 135.100 ;
        RECT 35.800 134.800 36.200 135.200 ;
        RECT 31.800 134.200 32.100 134.800 ;
        RECT 32.600 134.200 32.900 134.800 ;
        RECT 31.800 133.800 32.200 134.200 ;
        RECT 32.600 133.800 33.000 134.200 ;
        RECT 30.200 132.800 30.600 133.200 ;
        RECT 31.000 132.800 31.400 133.200 ;
        RECT 30.200 132.200 30.500 132.800 ;
        RECT 30.200 131.800 30.600 132.200 ;
        RECT 34.200 131.200 34.500 134.800 ;
        RECT 35.000 133.800 35.400 134.200 ;
        RECT 28.600 130.800 29.000 131.200 ;
        RECT 34.200 130.800 34.600 131.200 ;
        RECT 28.600 129.200 28.900 130.800 ;
        RECT 23.800 125.800 24.200 126.200 ;
        RECT 25.400 125.800 25.800 126.200 ;
        RECT 25.400 115.200 25.700 125.800 ;
        RECT 26.200 123.100 26.600 128.900 ;
        RECT 28.600 128.800 29.000 129.200 ;
        RECT 30.200 128.800 30.600 129.200 ;
        RECT 30.200 128.200 30.500 128.800 ;
        RECT 30.200 127.800 30.600 128.200 ;
        RECT 33.400 127.800 33.800 128.200 ;
        RECT 34.200 127.800 34.600 128.200 ;
        RECT 33.400 127.200 33.700 127.800 ;
        RECT 29.400 126.800 29.800 127.200 ;
        RECT 30.200 127.100 30.600 127.200 ;
        RECT 31.000 127.100 31.400 127.200 ;
        RECT 30.200 126.800 31.400 127.100 ;
        RECT 33.400 126.800 33.800 127.200 ;
        RECT 29.400 126.200 29.700 126.800 ;
        RECT 29.400 125.800 29.800 126.200 ;
        RECT 32.600 126.100 33.000 126.200 ;
        RECT 33.400 126.100 33.800 126.200 ;
        RECT 32.600 125.800 33.800 126.100 ;
        RECT 33.400 125.100 33.800 125.200 ;
        RECT 34.200 125.100 34.500 127.800 ;
        RECT 33.400 124.800 34.500 125.100 ;
        RECT 33.400 124.200 33.700 124.800 ;
        RECT 33.400 123.800 33.800 124.200 ;
        RECT 28.600 121.800 29.000 122.200 ;
        RECT 25.400 114.800 25.800 115.200 ;
        RECT 25.400 111.800 25.800 112.200 ;
        RECT 27.800 112.100 28.200 117.900 ;
        RECT 28.600 117.200 28.900 121.800 ;
        RECT 28.600 116.800 29.000 117.200 ;
        RECT 28.600 115.800 29.000 116.200 ;
        RECT 28.600 115.200 28.900 115.800 ;
        RECT 28.600 114.800 29.000 115.200 ;
        RECT 31.800 114.700 32.200 115.100 ;
        RECT 31.800 113.200 32.100 114.700 ;
        RECT 31.800 112.800 32.200 113.200 ;
        RECT 32.600 112.100 33.000 117.900 ;
        RECT 34.200 113.100 34.600 115.900 ;
        RECT 35.000 115.200 35.300 133.800 ;
        RECT 36.600 123.100 36.900 135.800 ;
        RECT 38.200 135.200 38.500 136.800 ;
        RECT 38.200 134.800 38.600 135.200 ;
        RECT 39.000 134.200 39.300 143.800 ;
        RECT 42.200 135.200 42.500 143.800 ;
        RECT 43.800 143.100 44.100 146.800 ;
        RECT 44.600 146.100 45.000 146.200 ;
        RECT 45.400 146.100 45.800 146.200 ;
        RECT 44.600 145.800 45.800 146.100 ;
        RECT 47.000 145.100 47.300 146.800 ;
        RECT 49.000 146.700 49.400 146.800 ;
        RECT 50.400 145.100 50.700 147.500 ;
        RECT 51.000 147.100 51.400 147.200 ;
        RECT 51.800 147.100 52.200 147.200 ;
        RECT 51.000 146.800 52.200 147.100 ;
        RECT 52.600 146.800 53.000 147.200 ;
        RECT 52.600 146.200 52.900 146.800 ;
        RECT 56.600 146.200 56.900 150.800 ;
        RECT 58.200 147.200 58.500 151.800 ;
        RECT 61.400 150.800 61.800 151.200 ;
        RECT 63.000 151.100 63.300 161.800 ;
        RECT 63.800 152.100 64.200 157.900 ;
        RECT 63.000 150.800 64.100 151.100 ;
        RECT 61.400 149.200 61.700 150.800 ;
        RECT 61.400 148.800 61.800 149.200 ;
        RECT 62.200 148.100 62.600 148.200 ;
        RECT 63.000 148.100 63.400 148.200 ;
        RECT 62.200 147.800 63.400 148.100 ;
        RECT 57.400 146.800 57.800 147.200 ;
        RECT 58.200 146.800 58.600 147.200 ;
        RECT 60.600 147.100 61.000 147.200 ;
        RECT 60.600 146.800 61.700 147.100 ;
        RECT 57.400 146.200 57.700 146.800 ;
        RECT 47.000 144.700 47.400 145.100 ;
        RECT 50.300 144.700 50.700 145.100 ;
        RECT 51.000 145.800 51.400 146.200 ;
        RECT 51.800 145.800 52.200 146.200 ;
        RECT 52.600 145.800 53.000 146.200 ;
        RECT 56.600 145.800 57.000 146.200 ;
        RECT 57.400 145.800 57.800 146.200 ;
        RECT 43.000 142.800 44.100 143.100 ;
        RECT 43.000 136.200 43.300 142.800 ;
        RECT 43.800 141.800 44.200 142.200 ;
        RECT 43.800 136.200 44.100 141.800 ;
        RECT 51.000 139.200 51.300 145.800 ;
        RECT 51.800 144.200 52.100 145.800 ;
        RECT 55.000 145.100 55.400 145.200 ;
        RECT 55.800 145.100 56.200 145.200 ;
        RECT 55.000 144.800 56.200 145.100 ;
        RECT 51.800 143.800 52.200 144.200 ;
        RECT 51.800 140.200 52.100 143.800 ;
        RECT 57.400 140.200 57.700 145.800 ;
        RECT 51.800 139.800 52.200 140.200 ;
        RECT 54.200 139.800 54.600 140.200 ;
        RECT 57.400 139.800 57.800 140.200 ;
        RECT 54.200 139.200 54.500 139.800 ;
        RECT 51.000 138.800 51.400 139.200 ;
        RECT 54.200 138.800 54.600 139.200 ;
        RECT 44.600 137.100 45.000 137.200 ;
        RECT 44.600 136.800 45.700 137.100 ;
        RECT 43.000 135.800 43.400 136.200 ;
        RECT 43.800 135.800 44.200 136.200 ;
        RECT 42.200 134.800 42.600 135.200 ;
        RECT 37.400 133.800 37.800 134.200 ;
        RECT 39.000 133.800 39.400 134.200 ;
        RECT 41.400 134.100 41.800 134.200 ;
        RECT 42.200 134.100 42.600 134.200 ;
        RECT 41.400 133.800 42.600 134.100 ;
        RECT 37.400 133.200 37.700 133.800 ;
        RECT 37.400 132.800 37.800 133.200 ;
        RECT 39.000 133.100 39.400 133.200 ;
        RECT 39.800 133.100 40.200 133.200 ;
        RECT 39.000 132.800 40.200 133.100 ;
        RECT 40.600 131.800 41.000 132.200 ;
        RECT 37.400 130.800 37.800 131.200 ;
        RECT 37.400 127.200 37.700 130.800 ;
        RECT 40.600 130.200 40.900 131.800 ;
        RECT 43.000 131.200 43.300 135.800 ;
        RECT 44.600 134.800 45.000 135.200 ;
        RECT 43.800 133.800 44.200 134.200 ;
        RECT 43.800 133.200 44.100 133.800 ;
        RECT 43.800 132.800 44.200 133.200 ;
        RECT 43.000 130.800 43.400 131.200 ;
        RECT 40.600 129.800 41.000 130.200 ;
        RECT 43.000 128.800 43.400 129.200 ;
        RECT 38.200 127.800 38.600 128.200 ;
        RECT 42.200 127.800 42.600 128.200 ;
        RECT 38.200 127.200 38.500 127.800 ;
        RECT 37.400 126.800 37.800 127.200 ;
        RECT 38.200 126.800 38.600 127.200 ;
        RECT 37.400 125.800 37.800 126.200 ;
        RECT 37.400 125.200 37.700 125.800 ;
        RECT 37.400 124.800 37.800 125.200 ;
        RECT 36.600 122.800 37.700 123.100 ;
        RECT 36.600 121.800 37.000 122.200 ;
        RECT 35.000 115.100 35.400 115.200 ;
        RECT 35.800 115.100 36.200 115.200 ;
        RECT 35.000 114.800 36.200 115.100 ;
        RECT 35.000 114.100 35.400 114.200 ;
        RECT 35.800 114.100 36.200 114.200 ;
        RECT 35.000 113.800 36.200 114.100 ;
        RECT 25.400 111.200 25.700 111.800 ;
        RECT 25.400 110.800 25.800 111.200 ;
        RECT 23.800 108.800 24.200 109.200 ;
        RECT 23.800 108.200 24.100 108.800 ;
        RECT 23.800 107.800 24.200 108.200 ;
        RECT 25.500 107.800 25.900 107.900 ;
        RECT 25.500 107.500 28.300 107.800 ;
        RECT 28.600 107.500 29.000 107.900 ;
        RECT 23.800 107.100 24.200 107.200 ;
        RECT 23.000 106.800 24.200 107.100 ;
        RECT 22.200 105.800 22.600 106.200 ;
        RECT 22.200 105.200 22.500 105.800 ;
        RECT 19.000 105.100 19.400 105.200 ;
        RECT 19.800 105.100 20.200 105.200 ;
        RECT 19.000 104.800 20.200 105.100 ;
        RECT 22.200 104.800 22.600 105.200 ;
        RECT 25.500 105.100 25.800 107.500 ;
        RECT 26.200 107.400 26.600 107.500 ;
        RECT 27.900 107.400 28.300 107.500 ;
        RECT 28.700 107.100 29.000 107.500 ;
        RECT 26.200 106.800 29.000 107.100 ;
        RECT 29.400 107.800 29.800 108.200 ;
        RECT 29.400 107.200 29.700 107.800 ;
        RECT 29.400 106.800 29.800 107.200 ;
        RECT 30.200 106.800 30.600 107.200 ;
        RECT 26.200 106.100 26.500 106.800 ;
        RECT 26.100 105.700 26.500 106.100 ;
        RECT 28.700 105.100 29.000 106.800 ;
        RECT 30.200 106.200 30.500 106.800 ;
        RECT 30.200 105.800 30.600 106.200 ;
        RECT 31.800 105.800 32.200 106.200 ;
        RECT 34.200 106.100 34.600 106.200 ;
        RECT 35.000 106.100 35.400 106.200 ;
        RECT 34.200 105.800 35.400 106.100 ;
        RECT 19.000 104.200 19.300 104.800 ;
        RECT 19.000 103.800 19.400 104.200 ;
        RECT 22.200 100.100 22.500 104.800 ;
        RECT 25.500 104.700 25.900 105.100 ;
        RECT 28.600 104.700 29.000 105.100 ;
        RECT 31.800 105.200 32.100 105.800 ;
        RECT 31.800 104.800 32.200 105.200 ;
        RECT 26.200 101.800 26.600 102.200 ;
        RECT 27.000 101.800 27.400 102.200 ;
        RECT 22.200 99.800 23.300 100.100 ;
        RECT 19.000 95.000 19.400 95.100 ;
        RECT 19.800 95.000 20.200 95.100 ;
        RECT 19.000 94.700 20.200 95.000 ;
        RECT 18.200 93.800 18.600 94.200 ;
        RECT 18.200 86.800 18.600 87.200 ;
        RECT 15.000 81.800 15.400 82.200 ;
        RECT 16.600 81.800 17.000 82.200 ;
        RECT 15.000 74.200 15.300 81.800 ;
        RECT 15.800 75.100 16.200 75.200 ;
        RECT 16.600 75.100 17.000 75.200 ;
        RECT 15.800 74.800 17.000 75.100 ;
        RECT 14.200 74.100 14.600 74.200 ;
        RECT 15.000 74.100 15.400 74.200 ;
        RECT 14.200 73.800 15.400 74.100 ;
        RECT 16.600 66.300 16.900 74.800 ;
        RECT 17.400 72.100 17.800 77.900 ;
        RECT 16.600 65.900 17.000 66.300 ;
        RECT 15.800 64.800 16.200 65.200 ;
        RECT 15.800 59.200 16.100 64.800 ;
        RECT 17.400 63.100 17.800 68.900 ;
        RECT 18.200 67.200 18.500 86.800 ;
        RECT 19.000 86.300 19.300 94.700 ;
        RECT 20.600 92.100 21.000 97.900 ;
        RECT 22.200 93.100 22.600 95.900 ;
        RECT 23.000 89.200 23.300 99.800 ;
        RECT 26.200 95.200 26.500 101.800 ;
        RECT 26.200 94.800 26.600 95.200 ;
        RECT 27.000 94.200 27.300 101.800 ;
        RECT 31.800 98.200 32.100 104.800 ;
        RECT 31.800 97.800 32.200 98.200 ;
        RECT 27.800 95.100 28.200 95.200 ;
        RECT 28.600 95.100 29.000 95.200 ;
        RECT 27.800 94.800 29.000 95.100 ;
        RECT 31.000 94.800 31.400 95.200 ;
        RECT 31.000 94.200 31.300 94.800 ;
        RECT 25.400 94.100 25.800 94.200 ;
        RECT 26.200 94.100 26.600 94.200 ;
        RECT 25.400 93.800 26.600 94.100 ;
        RECT 27.000 93.800 27.400 94.200 ;
        RECT 31.000 93.800 31.400 94.200 ;
        RECT 27.000 92.800 27.400 93.200 ;
        RECT 29.400 93.100 29.800 93.200 ;
        RECT 30.200 93.100 30.600 93.200 ;
        RECT 29.400 92.800 30.600 93.100 ;
        RECT 27.000 92.200 27.300 92.800 ;
        RECT 27.000 91.800 27.400 92.200 ;
        RECT 31.800 91.200 32.100 97.800 ;
        RECT 35.800 97.200 36.100 113.800 ;
        RECT 36.600 109.200 36.900 121.800 ;
        RECT 37.400 116.200 37.700 122.800 ;
        RECT 37.400 115.800 37.800 116.200 ;
        RECT 36.600 108.800 37.000 109.200 ;
        RECT 37.400 109.100 37.700 115.800 ;
        RECT 38.200 110.200 38.500 126.800 ;
        RECT 42.200 126.200 42.500 127.800 ;
        RECT 39.800 125.800 40.200 126.200 ;
        RECT 42.200 125.800 42.600 126.200 ;
        RECT 39.800 125.200 40.100 125.800 ;
        RECT 43.000 125.200 43.300 128.800 ;
        RECT 43.800 127.800 44.200 128.200 ;
        RECT 43.800 127.200 44.100 127.800 ;
        RECT 43.800 126.800 44.200 127.200 ;
        RECT 44.600 126.100 44.900 134.800 ;
        RECT 45.400 129.200 45.700 136.800 ;
        RECT 48.600 135.900 49.000 136.300 ;
        RECT 51.900 135.900 52.300 136.300 ;
        RECT 48.600 134.200 48.900 135.900 ;
        RECT 50.600 134.200 51.000 134.300 ;
        RECT 47.800 133.800 48.200 134.200 ;
        RECT 48.600 133.900 51.000 134.200 ;
        RECT 47.800 129.200 48.100 133.800 ;
        RECT 48.600 133.500 48.900 133.900 ;
        RECT 49.300 133.500 49.700 133.600 ;
        RECT 51.000 133.500 51.400 133.600 ;
        RECT 52.000 133.500 52.300 135.900 ;
        RECT 56.600 135.800 57.000 136.200 ;
        RECT 55.800 134.800 56.200 135.200 ;
        RECT 55.800 134.200 56.100 134.800 ;
        RECT 56.600 134.200 56.900 135.800 ;
        RECT 57.400 134.800 57.800 135.200 ;
        RECT 48.600 133.100 49.000 133.500 ;
        RECT 49.300 133.200 51.400 133.500 ;
        RECT 45.400 128.800 45.800 129.200 ;
        RECT 47.800 128.800 48.200 129.200 ;
        RECT 48.600 128.800 49.000 129.200 ;
        RECT 43.800 125.800 44.900 126.100 ;
        RECT 48.600 126.200 48.900 128.800 ;
        RECT 49.400 127.200 49.700 133.200 ;
        RECT 51.900 133.100 52.300 133.500 ;
        RECT 52.600 133.800 53.000 134.200 ;
        RECT 55.800 133.800 56.200 134.200 ;
        RECT 56.600 133.800 57.000 134.200 ;
        RECT 52.600 132.200 52.900 133.800 ;
        RECT 52.600 131.800 53.000 132.200 ;
        RECT 54.200 131.800 54.600 132.200 ;
        RECT 51.000 129.800 51.400 130.200 ;
        RECT 51.000 129.200 51.300 129.800 ;
        RECT 51.000 128.800 51.400 129.200 ;
        RECT 51.800 128.800 52.200 129.200 ;
        RECT 51.800 128.200 52.100 128.800 ;
        RECT 51.800 127.800 52.200 128.200 ;
        RECT 52.600 127.800 53.000 128.200 ;
        RECT 52.600 127.200 52.900 127.800 ;
        RECT 49.400 126.800 49.800 127.200 ;
        RECT 52.600 126.800 53.000 127.200 ;
        RECT 52.600 126.200 52.900 126.800 ;
        RECT 48.600 125.800 49.000 126.200 ;
        RECT 50.200 125.800 50.600 126.200 ;
        RECT 52.600 125.800 53.000 126.200 ;
        RECT 39.800 124.800 40.200 125.200 ;
        RECT 42.200 124.800 42.600 125.200 ;
        RECT 43.000 124.800 43.400 125.200 ;
        RECT 39.000 124.100 39.400 124.200 ;
        RECT 39.800 124.100 40.200 124.200 ;
        RECT 39.000 123.800 40.200 124.100 ;
        RECT 40.600 124.100 41.000 124.200 ;
        RECT 41.400 124.100 41.800 124.200 ;
        RECT 40.600 123.800 41.800 124.100 ;
        RECT 42.200 123.200 42.500 124.800 ;
        RECT 42.200 122.800 42.600 123.200 ;
        RECT 43.800 119.200 44.100 125.800 ;
        RECT 50.200 125.200 50.500 125.800 ;
        RECT 50.200 124.800 50.600 125.200 ;
        RECT 50.200 121.800 50.600 122.200 ;
        RECT 47.800 119.800 48.200 120.200 ;
        RECT 43.800 118.800 44.200 119.200 ;
        RECT 39.800 117.800 40.200 118.200 ;
        RECT 39.800 114.200 40.100 117.800 ;
        RECT 42.200 117.100 42.600 117.200 ;
        RECT 43.000 117.100 43.400 117.200 ;
        RECT 42.200 116.800 43.400 117.100 ;
        RECT 43.800 117.100 44.200 117.200 ;
        RECT 44.600 117.100 45.000 117.200 ;
        RECT 43.800 116.800 45.000 117.100 ;
        RECT 47.800 116.200 48.100 119.800 ;
        RECT 48.600 117.100 49.000 117.200 ;
        RECT 49.400 117.100 49.800 117.200 ;
        RECT 48.600 116.800 49.800 117.100 ;
        RECT 50.200 116.200 50.500 121.800 ;
        RECT 51.800 118.800 52.200 119.200 ;
        RECT 51.800 118.200 52.100 118.800 ;
        RECT 51.800 117.800 52.200 118.200 ;
        RECT 51.000 117.100 51.400 117.200 ;
        RECT 51.800 117.100 52.200 117.200 ;
        RECT 52.600 117.100 53.000 117.200 ;
        RECT 51.000 116.800 53.000 117.100 ;
        RECT 54.200 116.200 54.500 131.800 ;
        RECT 56.600 130.800 57.000 131.200 ;
        RECT 55.000 126.100 55.400 126.200 ;
        RECT 55.800 126.100 56.200 126.200 ;
        RECT 55.000 125.800 56.200 126.100 ;
        RECT 55.800 124.800 56.200 125.200 ;
        RECT 55.800 124.200 56.100 124.800 ;
        RECT 55.800 123.800 56.200 124.200 ;
        RECT 55.000 121.800 55.400 122.200 ;
        RECT 55.000 121.200 55.300 121.800 ;
        RECT 55.000 120.800 55.400 121.200 ;
        RECT 56.600 120.200 56.900 130.800 ;
        RECT 57.400 130.200 57.700 134.800 ;
        RECT 57.400 129.800 57.800 130.200 ;
        RECT 58.200 129.100 58.500 146.800 ;
        RECT 59.000 146.100 59.400 146.200 ;
        RECT 59.800 146.100 60.200 146.200 ;
        RECT 59.000 145.800 60.200 146.100 ;
        RECT 59.000 141.800 59.400 142.200 ;
        RECT 59.000 136.200 59.300 141.800 ;
        RECT 61.400 139.200 61.700 146.800 ;
        RECT 63.800 146.200 64.100 150.800 ;
        RECT 64.600 149.200 64.900 163.800 ;
        RECT 65.400 163.100 65.800 168.900 ;
        RECT 69.400 166.800 69.800 167.200 ;
        RECT 66.200 166.100 66.600 166.200 ;
        RECT 67.000 166.100 67.400 166.200 ;
        RECT 66.200 165.800 67.400 166.100 ;
        RECT 67.000 154.800 67.400 155.200 ;
        RECT 67.000 151.200 67.300 154.800 ;
        RECT 68.600 152.100 69.000 157.900 ;
        RECT 69.400 154.200 69.700 166.800 ;
        RECT 70.200 163.100 70.600 168.900 ;
        RECT 71.800 165.100 72.200 167.900 ;
        RECT 72.600 164.800 73.000 165.200 ;
        RECT 72.600 162.200 72.900 164.800 ;
        RECT 75.000 163.100 75.400 168.900 ;
        RECT 79.000 165.900 79.400 166.300 ;
        RECT 72.600 161.800 73.000 162.200 ;
        RECT 72.600 156.200 72.900 161.800 ;
        RECT 69.400 153.800 69.800 154.200 ;
        RECT 69.400 153.200 69.700 153.800 ;
        RECT 69.400 152.800 69.800 153.200 ;
        RECT 70.200 153.100 70.600 155.900 ;
        RECT 72.600 155.800 73.000 156.200 ;
        RECT 71.000 151.800 71.400 152.200 ;
        RECT 71.000 151.200 71.300 151.800 ;
        RECT 67.000 150.800 67.400 151.200 ;
        RECT 71.000 150.800 71.400 151.200 ;
        RECT 68.600 149.800 69.000 150.200 ;
        RECT 68.600 149.200 68.900 149.800 ;
        RECT 64.600 148.800 65.000 149.200 ;
        RECT 68.600 148.800 69.000 149.200 ;
        RECT 71.000 148.800 71.400 149.200 ;
        RECT 71.000 148.200 71.300 148.800 ;
        RECT 71.000 147.800 71.400 148.200 ;
        RECT 67.000 146.800 67.400 147.200 ;
        RECT 63.000 145.800 63.400 146.200 ;
        RECT 63.800 145.800 64.200 146.200 ;
        RECT 66.200 145.800 66.600 146.200 ;
        RECT 63.000 144.200 63.300 145.800 ;
        RECT 63.000 143.800 63.400 144.200 ;
        RECT 63.000 139.200 63.300 143.800 ;
        RECT 63.800 143.200 64.100 145.800 ;
        RECT 63.800 142.800 64.200 143.200 ;
        RECT 66.200 141.200 66.500 145.800 ;
        RECT 66.200 140.800 66.600 141.200 ;
        RECT 67.000 139.200 67.300 146.800 ;
        RECT 72.600 146.200 72.900 155.800 ;
        RECT 73.400 152.100 73.800 157.900 ;
        RECT 77.400 154.700 77.800 155.100 ;
        RECT 77.400 154.200 77.700 154.700 ;
        RECT 77.400 153.800 77.800 154.200 ;
        RECT 77.400 152.800 77.800 153.200 ;
        RECT 73.400 146.800 73.800 147.200 ;
        RECT 70.200 145.800 70.600 146.200 ;
        RECT 72.600 145.800 73.000 146.200 ;
        RECT 61.400 138.800 61.800 139.200 ;
        RECT 63.000 138.800 63.400 139.200 ;
        RECT 67.000 138.800 67.400 139.200 ;
        RECT 70.200 138.200 70.500 145.800 ;
        RECT 71.000 145.100 71.400 145.200 ;
        RECT 71.800 145.100 72.200 145.200 ;
        RECT 71.000 144.800 72.200 145.100 ;
        RECT 73.400 143.200 73.700 146.800 ;
        RECT 73.400 142.800 73.800 143.200 ;
        RECT 76.600 143.100 77.000 148.900 ;
        RECT 77.400 147.200 77.700 152.800 ;
        RECT 78.200 152.100 78.600 157.900 ;
        RECT 77.400 146.800 77.800 147.200 ;
        RECT 78.200 146.800 78.600 147.200 ;
        RECT 74.200 142.100 74.600 142.200 ;
        RECT 75.000 142.100 75.400 142.200 ;
        RECT 74.200 141.800 75.400 142.100 ;
        RECT 78.200 139.200 78.500 146.800 ;
        RECT 79.000 146.100 79.300 165.900 ;
        RECT 79.800 163.100 80.200 168.900 ;
        RECT 80.600 166.800 81.000 167.200 ;
        RECT 80.600 163.200 80.900 166.800 ;
        RECT 81.400 165.100 81.800 167.900 ;
        RECT 84.600 167.800 85.000 168.200 ;
        RECT 90.200 167.800 90.600 168.200 ;
        RECT 80.600 162.800 81.000 163.200 ;
        RECT 82.200 162.800 82.600 163.200 ;
        RECT 82.200 157.200 82.500 162.800 ;
        RECT 82.200 156.800 82.600 157.200 ;
        RECT 79.800 153.100 80.200 155.900 ;
        RECT 80.600 151.800 81.000 152.200 ;
        RECT 83.000 152.100 83.400 157.900 ;
        RECT 84.600 154.200 84.900 167.800 ;
        RECT 86.200 166.100 86.600 166.200 ;
        RECT 87.000 166.100 87.400 166.200 ;
        RECT 86.200 165.800 87.400 166.100 ;
        RECT 88.600 166.100 89.000 166.200 ;
        RECT 89.400 166.100 89.800 166.200 ;
        RECT 88.600 165.800 89.800 166.100 ;
        RECT 87.000 154.700 87.400 155.200 ;
        RECT 84.600 153.800 85.000 154.200 ;
        RECT 80.600 151.200 80.900 151.800 ;
        RECT 80.600 150.800 81.000 151.200 ;
        RECT 87.000 151.100 87.300 154.700 ;
        RECT 87.800 152.100 88.200 157.900 ;
        RECT 88.600 153.800 89.000 154.200 ;
        RECT 87.000 150.800 88.100 151.100 ;
        RECT 87.800 149.200 88.100 150.800 ;
        RECT 79.800 146.200 80.200 146.300 ;
        RECT 80.600 146.200 81.000 146.300 ;
        RECT 79.800 146.100 81.000 146.200 ;
        RECT 79.000 145.900 81.000 146.100 ;
        RECT 79.000 145.800 80.100 145.900 ;
        RECT 80.600 143.800 81.000 144.200 ;
        RECT 78.200 138.800 78.600 139.200 ;
        RECT 63.800 137.800 64.200 138.200 ;
        RECT 70.200 137.800 70.600 138.200 ;
        RECT 63.800 136.200 64.100 137.800 ;
        RECT 64.600 137.100 65.000 137.200 ;
        RECT 66.200 137.100 66.600 137.200 ;
        RECT 64.600 136.800 66.600 137.100 ;
        RECT 67.800 137.100 68.200 137.200 ;
        RECT 67.800 136.800 68.900 137.100 ;
        RECT 66.200 136.200 66.500 136.800 ;
        RECT 59.000 135.800 59.400 136.200 ;
        RECT 61.400 135.800 61.800 136.200 ;
        RECT 63.000 135.800 63.400 136.200 ;
        RECT 63.800 135.800 64.200 136.200 ;
        RECT 66.200 135.800 66.600 136.200 ;
        RECT 59.000 134.200 59.300 135.800 ;
        RECT 61.400 135.200 61.700 135.800 ;
        RECT 63.000 135.200 63.300 135.800 ;
        RECT 61.400 134.800 61.800 135.200 ;
        RECT 63.000 134.800 63.400 135.200 ;
        RECT 63.800 134.800 64.200 135.200 ;
        RECT 59.000 133.800 59.400 134.200 ;
        RECT 61.400 134.100 61.800 134.200 ;
        RECT 62.200 134.100 62.600 134.200 ;
        RECT 61.400 133.800 62.600 134.100 ;
        RECT 57.400 128.800 58.500 129.100 ;
        RECT 57.400 128.200 57.700 128.800 ;
        RECT 57.400 127.800 57.800 128.200 ;
        RECT 59.000 128.100 59.400 128.200 ;
        RECT 59.800 128.100 60.200 128.200 ;
        RECT 59.000 127.800 60.200 128.100 ;
        RECT 56.600 119.800 57.000 120.200 ;
        RECT 56.600 116.200 56.900 119.800 ;
        RECT 45.400 115.800 45.800 116.200 ;
        RECT 47.800 115.800 48.200 116.200 ;
        RECT 50.200 115.800 50.600 116.200 ;
        RECT 51.000 115.800 51.400 116.200 ;
        RECT 54.200 115.800 54.600 116.200 ;
        RECT 55.000 116.100 55.400 116.200 ;
        RECT 55.800 116.100 56.200 116.200 ;
        RECT 55.000 115.800 56.200 116.100 ;
        RECT 56.600 115.800 57.000 116.200 ;
        RECT 45.400 115.200 45.700 115.800 ;
        RECT 40.600 114.800 41.000 115.200 ;
        RECT 43.000 114.800 43.400 115.200 ;
        RECT 45.400 114.800 45.800 115.200 ;
        RECT 49.400 115.100 49.800 115.200 ;
        RECT 50.200 115.100 50.600 115.200 ;
        RECT 49.400 114.800 50.600 115.100 ;
        RECT 40.600 114.200 40.900 114.800 ;
        RECT 39.800 113.800 40.200 114.200 ;
        RECT 40.600 113.800 41.000 114.200 ;
        RECT 39.000 112.800 39.400 113.200 ;
        RECT 41.400 112.800 41.800 113.200 ;
        RECT 39.000 112.200 39.300 112.800 ;
        RECT 39.000 111.800 39.400 112.200 ;
        RECT 38.200 109.800 38.600 110.200 ;
        RECT 39.800 109.800 40.200 110.200 ;
        RECT 37.400 108.800 38.500 109.100 ;
        RECT 36.600 108.100 37.000 108.200 ;
        RECT 37.400 108.100 37.800 108.200 ;
        RECT 36.600 107.800 37.800 108.100 ;
        RECT 36.600 107.100 37.000 107.200 ;
        RECT 37.400 107.100 37.800 107.200 ;
        RECT 36.600 106.800 37.800 107.100 ;
        RECT 37.400 103.800 37.800 104.200 ;
        RECT 35.000 96.800 35.400 97.200 ;
        RECT 35.800 96.800 36.200 97.200 ;
        RECT 35.000 96.200 35.300 96.800 ;
        RECT 33.400 95.800 33.800 96.200 ;
        RECT 35.000 95.800 35.400 96.200 ;
        RECT 33.400 95.200 33.700 95.800 ;
        RECT 33.400 94.800 33.800 95.200 ;
        RECT 35.800 94.200 36.100 96.800 ;
        RECT 37.400 95.200 37.700 103.800 ;
        RECT 38.200 96.200 38.500 108.800 ;
        RECT 39.800 105.200 40.100 109.800 ;
        RECT 40.600 107.800 41.000 108.200 ;
        RECT 40.600 106.200 40.900 107.800 ;
        RECT 41.400 107.200 41.700 112.800 ;
        RECT 43.000 108.200 43.300 114.800 ;
        RECT 51.000 114.200 51.300 115.800 ;
        RECT 53.400 115.100 53.800 115.200 ;
        RECT 54.200 115.100 54.600 115.200 ;
        RECT 53.400 114.800 54.600 115.100 ;
        RECT 51.000 113.800 51.400 114.200 ;
        RECT 57.400 114.100 57.700 127.800 ;
        RECT 61.400 127.200 61.700 133.800 ;
        RECT 63.800 131.200 64.100 134.800 ;
        RECT 65.400 133.800 65.800 134.200 ;
        RECT 65.400 132.200 65.700 133.800 ;
        RECT 65.400 131.800 65.800 132.200 ;
        RECT 63.800 130.800 64.200 131.200 ;
        RECT 65.400 129.200 65.700 131.800 ;
        RECT 65.400 128.800 65.800 129.200 ;
        RECT 66.200 128.100 66.500 135.800 ;
        RECT 67.000 135.100 67.400 135.200 ;
        RECT 67.800 135.100 68.200 135.200 ;
        RECT 67.000 134.800 68.200 135.100 ;
        RECT 68.600 132.200 68.900 136.800 ;
        RECT 71.000 136.800 71.400 137.200 ;
        RECT 71.800 136.800 72.200 137.200 ;
        RECT 73.400 137.100 73.800 137.200 ;
        RECT 74.200 137.100 74.600 137.200 ;
        RECT 73.400 136.800 74.600 137.100 ;
        RECT 71.000 136.200 71.300 136.800 ;
        RECT 71.800 136.200 72.100 136.800 ;
        RECT 71.000 135.800 71.400 136.200 ;
        RECT 71.800 135.800 72.200 136.200 ;
        RECT 75.700 135.900 76.100 136.300 ;
        RECT 79.000 135.900 79.400 136.300 ;
        RECT 71.000 135.200 71.300 135.800 ;
        RECT 69.400 134.800 69.800 135.200 ;
        RECT 71.000 134.800 71.400 135.200 ;
        RECT 72.600 134.800 73.000 135.200 ;
        RECT 69.400 134.200 69.700 134.800 ;
        RECT 72.600 134.200 72.900 134.800 ;
        RECT 69.400 133.800 69.800 134.200 ;
        RECT 71.000 133.800 71.400 134.200 ;
        RECT 72.600 133.800 73.000 134.200 ;
        RECT 73.400 134.100 73.800 134.200 ;
        RECT 74.200 134.100 74.600 134.200 ;
        RECT 73.400 133.800 74.600 134.100 ;
        RECT 75.000 133.800 75.400 134.200 ;
        RECT 68.600 131.800 69.000 132.200 ;
        RECT 65.400 127.800 66.500 128.100 ;
        RECT 61.400 126.800 61.800 127.200 ;
        RECT 63.800 126.800 64.200 127.200 ;
        RECT 61.400 125.200 61.700 126.800 ;
        RECT 63.000 125.800 63.400 126.200 ;
        RECT 63.000 125.200 63.300 125.800 ;
        RECT 59.800 124.800 60.200 125.200 ;
        RECT 61.400 124.800 61.800 125.200 ;
        RECT 63.000 124.800 63.400 125.200 ;
        RECT 58.200 124.100 58.600 124.200 ;
        RECT 59.000 124.100 59.400 124.200 ;
        RECT 58.200 123.800 59.400 124.100 ;
        RECT 59.800 116.200 60.100 124.800 ;
        RECT 59.000 116.100 59.400 116.200 ;
        RECT 59.800 116.100 60.200 116.200 ;
        RECT 59.000 115.800 60.200 116.100 ;
        RECT 62.200 116.100 62.600 116.200 ;
        RECT 63.000 116.100 63.400 116.200 ;
        RECT 62.200 115.800 63.400 116.100 ;
        RECT 58.200 115.100 58.600 115.200 ;
        RECT 59.000 115.100 59.400 115.200 ;
        RECT 58.200 114.800 59.400 115.100 ;
        RECT 60.600 114.800 61.000 115.200 ;
        RECT 61.400 114.800 61.800 115.200 ;
        RECT 58.200 114.100 58.600 114.200 ;
        RECT 57.400 113.800 58.600 114.100 ;
        RECT 51.000 111.200 51.300 113.800 ;
        RECT 56.600 113.100 57.000 113.200 ;
        RECT 57.400 113.100 57.800 113.200 ;
        RECT 56.600 112.800 57.800 113.100 ;
        RECT 57.400 111.800 57.800 112.200 ;
        RECT 51.000 110.800 51.400 111.200 ;
        RECT 46.200 108.800 46.600 109.200 ;
        RECT 43.000 107.800 43.400 108.200 ;
        RECT 44.600 107.800 45.000 108.200 ;
        RECT 41.400 106.800 41.800 107.200 ;
        RECT 43.000 106.800 43.400 107.200 ;
        RECT 40.600 105.800 41.000 106.200 ;
        RECT 39.000 104.800 39.400 105.200 ;
        RECT 39.800 104.800 40.200 105.200 ;
        RECT 40.600 104.800 41.000 105.200 ;
        RECT 39.000 104.200 39.300 104.800 ;
        RECT 39.000 103.800 39.400 104.200 ;
        RECT 39.800 99.200 40.100 104.800 ;
        RECT 40.600 103.200 40.900 104.800 ;
        RECT 41.400 104.100 41.800 104.200 ;
        RECT 42.200 104.100 42.600 104.200 ;
        RECT 41.400 103.800 42.600 104.100 ;
        RECT 40.600 102.800 41.000 103.200 ;
        RECT 39.800 98.800 40.200 99.200 ;
        RECT 38.200 95.800 38.600 96.200 ;
        RECT 41.400 95.800 41.800 96.200 ;
        RECT 36.600 94.800 37.000 95.200 ;
        RECT 37.400 94.800 37.800 95.200 ;
        RECT 38.200 94.800 38.600 95.200 ;
        RECT 39.000 95.100 39.400 95.200 ;
        RECT 39.800 95.100 40.200 95.200 ;
        RECT 39.000 94.800 40.200 95.100 ;
        RECT 32.600 94.100 33.000 94.200 ;
        RECT 33.400 94.100 33.800 94.200 ;
        RECT 32.600 93.800 33.800 94.100 ;
        RECT 34.200 93.800 34.600 94.200 ;
        RECT 35.800 93.800 36.200 94.200 ;
        RECT 34.200 93.200 34.500 93.800 ;
        RECT 34.200 92.800 34.600 93.200 ;
        RECT 34.200 91.800 34.600 92.200 ;
        RECT 27.000 90.800 27.400 91.200 ;
        RECT 31.800 90.800 32.200 91.200 ;
        RECT 27.000 89.200 27.300 90.800 ;
        RECT 34.200 89.200 34.500 91.800 ;
        RECT 36.600 90.200 36.900 94.800 ;
        RECT 38.200 94.200 38.500 94.800 ;
        RECT 41.400 94.200 41.700 95.800 ;
        RECT 43.000 95.100 43.300 106.800 ;
        RECT 44.600 97.200 44.900 107.800 ;
        RECT 46.200 104.200 46.500 108.800 ;
        RECT 55.000 106.800 55.400 107.200 ;
        RECT 55.000 106.200 55.300 106.800 ;
        RECT 57.400 106.200 57.700 111.800 ;
        RECT 47.000 106.100 47.400 106.200 ;
        RECT 47.800 106.100 48.200 106.200 ;
        RECT 47.000 105.800 48.200 106.100 ;
        RECT 53.400 105.800 53.800 106.200 ;
        RECT 54.200 105.800 54.600 106.200 ;
        RECT 55.000 105.800 55.400 106.200 ;
        RECT 57.400 105.800 57.800 106.200 ;
        RECT 46.200 103.800 46.600 104.200 ;
        RECT 53.400 102.200 53.700 105.800 ;
        RECT 51.800 101.800 52.200 102.200 ;
        RECT 53.400 101.800 53.800 102.200 ;
        RECT 44.600 96.800 45.000 97.200 ;
        RECT 49.400 95.900 49.800 96.300 ;
        RECT 42.200 94.800 43.300 95.100 ;
        RECT 46.200 95.100 46.600 95.200 ;
        RECT 47.000 95.100 47.400 95.200 ;
        RECT 46.200 94.800 47.400 95.100 ;
        RECT 47.800 94.800 48.200 95.200 ;
        RECT 38.200 93.800 38.600 94.200 ;
        RECT 39.000 93.800 39.400 94.200 ;
        RECT 39.800 93.800 40.200 94.200 ;
        RECT 41.400 93.800 41.800 94.200 ;
        RECT 39.000 93.200 39.300 93.800 ;
        RECT 39.000 92.800 39.400 93.200 ;
        RECT 36.600 89.800 37.000 90.200 ;
        RECT 39.800 89.200 40.100 93.800 ;
        RECT 42.200 92.200 42.500 94.800 ;
        RECT 47.800 94.200 48.100 94.800 ;
        RECT 49.400 94.200 49.700 95.900 ;
        RECT 51.800 95.200 52.100 101.800 ;
        RECT 54.200 101.200 54.500 105.800 ;
        RECT 55.800 101.800 56.200 102.200 ;
        RECT 54.200 100.800 54.600 101.200 ;
        RECT 54.200 97.800 54.600 98.200 ;
        RECT 53.400 96.800 53.800 97.200 ;
        RECT 52.700 95.900 53.100 96.300 ;
        RECT 51.800 94.800 52.200 95.200 ;
        RECT 51.400 94.200 51.800 94.300 ;
        RECT 43.000 94.100 43.400 94.200 ;
        RECT 43.800 94.100 44.200 94.200 ;
        RECT 43.000 93.800 44.200 94.100 ;
        RECT 46.200 93.800 46.600 94.200 ;
        RECT 47.000 93.800 47.400 94.200 ;
        RECT 47.800 93.800 48.200 94.200 ;
        RECT 49.400 93.900 51.800 94.200 ;
        RECT 46.200 93.200 46.500 93.800 ;
        RECT 43.000 93.100 43.400 93.200 ;
        RECT 43.800 93.100 44.200 93.200 ;
        RECT 43.000 92.800 44.200 93.100 ;
        RECT 46.200 92.800 46.600 93.200 ;
        RECT 42.200 91.800 42.600 92.200 ;
        RECT 44.600 91.800 45.000 92.200 ;
        RECT 40.600 89.800 41.000 90.200 ;
        RECT 19.000 85.900 19.400 86.300 ;
        RECT 19.800 83.100 20.200 88.900 ;
        RECT 23.000 88.800 23.400 89.200 ;
        RECT 27.000 88.800 27.400 89.200 ;
        RECT 34.200 88.800 34.600 89.200 ;
        RECT 39.800 88.800 40.200 89.200 ;
        RECT 31.800 88.100 32.200 88.200 ;
        RECT 32.600 88.100 33.000 88.200 ;
        RECT 21.400 85.100 21.800 87.900 ;
        RECT 31.800 87.800 33.000 88.100 ;
        RECT 35.000 87.800 35.400 88.200 ;
        RECT 38.200 87.800 38.600 88.200 ;
        RECT 23.800 86.800 24.200 87.200 ;
        RECT 27.800 87.100 28.200 87.200 ;
        RECT 28.600 87.100 29.000 87.200 ;
        RECT 27.800 86.800 29.000 87.100 ;
        RECT 30.200 86.800 30.600 87.200 ;
        RECT 19.000 73.100 19.400 75.900 ;
        RECT 19.800 73.100 20.200 75.900 ;
        RECT 21.400 72.100 21.800 77.900 ;
        RECT 23.000 74.800 23.400 75.200 ;
        RECT 23.000 72.200 23.300 74.800 ;
        RECT 23.000 71.800 23.400 72.200 ;
        RECT 23.800 68.200 24.100 86.800 ;
        RECT 30.200 86.200 30.500 86.800 ;
        RECT 25.400 85.800 25.800 86.200 ;
        RECT 30.200 85.800 30.600 86.200 ;
        RECT 25.400 83.200 25.700 85.800 ;
        RECT 25.400 82.800 25.800 83.200 ;
        RECT 18.200 66.800 18.600 67.200 ;
        RECT 18.200 66.200 18.500 66.800 ;
        RECT 18.200 65.800 18.600 66.200 ;
        RECT 19.000 65.100 19.400 67.900 ;
        RECT 23.800 67.800 24.200 68.200 ;
        RECT 22.200 65.800 22.600 66.200 ;
        RECT 19.800 64.800 20.200 65.200 ;
        RECT 19.800 64.200 20.100 64.800 ;
        RECT 19.800 63.800 20.200 64.200 ;
        RECT 22.200 62.200 22.500 65.800 ;
        RECT 24.600 65.100 25.000 67.900 ;
        RECT 18.200 61.800 18.600 62.200 ;
        RECT 22.200 61.800 22.600 62.200 ;
        RECT 18.200 59.200 18.500 61.800 ;
        RECT 15.800 58.800 16.200 59.200 ;
        RECT 18.200 58.800 18.600 59.200 ;
        RECT 25.400 57.200 25.700 82.800 ;
        RECT 28.600 81.800 29.000 82.200 ;
        RECT 28.600 79.200 28.900 81.800 ;
        RECT 31.800 79.200 32.100 87.800 ;
        RECT 35.000 87.200 35.300 87.800 ;
        RECT 38.200 87.200 38.500 87.800 ;
        RECT 35.000 86.800 35.400 87.200 ;
        RECT 35.800 87.100 36.200 87.200 ;
        RECT 36.600 87.100 37.000 87.200 ;
        RECT 35.800 86.800 37.000 87.100 ;
        RECT 38.200 86.800 38.600 87.200 ;
        RECT 39.000 86.800 39.400 87.200 ;
        RECT 34.200 84.800 34.600 85.200 ;
        RECT 35.000 85.100 35.400 85.200 ;
        RECT 35.800 85.100 36.200 85.200 ;
        RECT 35.000 84.800 36.200 85.100 ;
        RECT 33.400 81.800 33.800 82.200 ;
        RECT 28.600 78.800 29.000 79.200 ;
        RECT 31.800 78.800 32.200 79.200 ;
        RECT 26.200 72.100 26.600 77.900 ;
        RECT 31.800 77.200 32.100 78.800 ;
        RECT 31.800 76.800 32.200 77.200 ;
        RECT 31.000 75.800 31.400 76.200 ;
        RECT 31.000 75.200 31.300 75.800 ;
        RECT 31.000 74.800 31.400 75.200 ;
        RECT 28.600 73.100 29.000 73.200 ;
        RECT 29.400 73.100 29.800 73.200 ;
        RECT 28.600 72.800 29.800 73.100 ;
        RECT 30.200 71.800 30.600 72.200 ;
        RECT 31.800 71.800 32.200 72.200 ;
        RECT 26.200 63.100 26.600 68.900 ;
        RECT 27.000 66.800 27.400 67.200 ;
        RECT 19.800 56.800 20.200 57.200 ;
        RECT 25.400 56.800 25.800 57.200 ;
        RECT 16.600 55.800 17.000 56.200 ;
        RECT 13.400 54.800 13.800 55.200 ;
        RECT 16.600 54.200 16.900 55.800 ;
        RECT 19.800 55.200 20.100 56.800 ;
        RECT 23.000 55.800 23.400 56.200 ;
        RECT 23.000 55.200 23.300 55.800 ;
        RECT 19.800 54.800 20.200 55.200 ;
        RECT 22.200 54.800 22.600 55.200 ;
        RECT 23.000 54.800 23.400 55.200 ;
        RECT 23.800 54.800 24.200 55.200 ;
        RECT 22.200 54.200 22.500 54.800 ;
        RECT 14.200 54.100 14.600 54.200 ;
        RECT 15.000 54.100 15.400 54.200 ;
        RECT 14.200 53.800 15.400 54.100 ;
        RECT 16.600 53.800 17.000 54.200 ;
        RECT 22.200 53.800 22.600 54.200 ;
        RECT 23.800 53.200 24.100 54.800 ;
        RECT 24.600 53.800 25.000 54.200 ;
        RECT 24.600 53.200 24.900 53.800 ;
        RECT 20.600 52.800 21.000 53.200 ;
        RECT 23.800 52.800 24.200 53.200 ;
        RECT 24.600 52.800 25.000 53.200 ;
        RECT 18.200 49.800 18.600 50.200 ;
        RECT 11.800 48.800 12.900 49.100 ;
        RECT 11.800 45.100 12.200 47.900 ;
        RECT 12.600 46.200 12.900 48.800 ;
        RECT 13.400 48.100 13.800 48.200 ;
        RECT 14.200 48.100 14.600 48.200 ;
        RECT 13.400 47.800 14.600 48.100 ;
        RECT 12.600 45.800 13.000 46.200 ;
        RECT 14.200 45.800 14.600 46.200 ;
        RECT 9.400 39.800 9.800 40.200 ;
        RECT 9.400 39.100 9.800 39.200 ;
        RECT 10.200 39.100 10.600 39.200 ;
        RECT 9.400 38.800 10.600 39.100 ;
        RECT 8.600 33.800 9.000 34.200 ;
        RECT 6.200 29.800 6.600 30.200 ;
        RECT 8.600 29.100 8.900 33.800 ;
        RECT 9.400 33.100 9.800 35.900 ;
        RECT 12.600 32.100 13.000 37.900 ;
        RECT 14.200 35.200 14.500 45.800 ;
        RECT 15.000 45.100 15.400 47.900 ;
        RECT 15.800 47.800 16.200 48.200 ;
        RECT 15.800 47.200 16.100 47.800 ;
        RECT 15.800 46.800 16.200 47.200 ;
        RECT 16.600 43.100 17.000 48.900 ;
        RECT 18.200 46.200 18.500 49.800 ;
        RECT 20.600 47.200 20.900 52.800 ;
        RECT 21.400 51.800 21.800 52.200 ;
        RECT 21.400 50.200 21.700 51.800 ;
        RECT 21.400 49.800 21.800 50.200 ;
        RECT 23.800 49.200 24.100 52.800 ;
        RECT 20.600 46.800 21.000 47.200 ;
        RECT 18.200 45.800 18.600 46.200 ;
        RECT 21.400 43.100 21.800 48.900 ;
        RECT 23.800 48.800 24.200 49.200 ;
        RECT 24.600 45.100 25.000 47.900 ;
        RECT 26.200 43.100 26.600 48.900 ;
        RECT 27.000 48.200 27.300 66.800 ;
        RECT 29.400 66.100 29.800 66.200 ;
        RECT 30.200 66.100 30.500 71.800 ;
        RECT 29.400 65.800 30.500 66.100 ;
        RECT 28.600 64.800 29.000 65.200 ;
        RECT 27.800 63.800 28.200 64.200 ;
        RECT 27.800 55.200 28.100 63.800 ;
        RECT 28.600 59.200 28.900 64.800 ;
        RECT 31.000 63.100 31.400 68.900 ;
        RECT 29.400 61.800 29.800 62.200 ;
        RECT 28.600 58.800 29.000 59.200 ;
        RECT 29.400 56.200 29.700 61.800 ;
        RECT 29.400 55.800 29.800 56.200 ;
        RECT 31.100 55.900 31.500 56.300 ;
        RECT 31.800 56.200 32.100 71.800 ;
        RECT 33.400 69.200 33.700 81.800 ;
        RECT 34.200 81.200 34.500 84.800 ;
        RECT 34.200 80.800 34.600 81.200 ;
        RECT 34.200 72.100 34.600 77.900 ;
        RECT 36.600 74.200 36.900 86.800 ;
        RECT 37.400 85.100 37.800 85.200 ;
        RECT 38.200 85.100 38.600 85.200 ;
        RECT 37.400 84.800 38.600 85.100 ;
        RECT 39.000 79.200 39.300 86.800 ;
        RECT 40.600 85.200 40.900 89.800 ;
        RECT 44.600 89.200 44.900 91.800 ;
        RECT 44.600 88.800 45.000 89.200 ;
        RECT 45.400 88.800 45.800 89.200 ;
        RECT 45.400 88.200 45.700 88.800 ;
        RECT 43.800 88.100 44.200 88.200 ;
        RECT 44.600 88.100 45.000 88.200 ;
        RECT 43.800 87.800 45.000 88.100 ;
        RECT 45.400 87.800 45.800 88.200 ;
        RECT 43.800 87.100 44.200 87.200 ;
        RECT 44.600 87.100 45.000 87.200 ;
        RECT 43.800 86.800 45.000 87.100 ;
        RECT 47.000 86.200 47.300 93.800 ;
        RECT 49.400 93.500 49.700 93.900 ;
        RECT 50.100 93.500 50.500 93.600 ;
        RECT 51.800 93.500 52.200 93.600 ;
        RECT 52.800 93.500 53.100 95.900 ;
        RECT 53.400 94.200 53.700 96.800 ;
        RECT 54.200 96.200 54.500 97.800 ;
        RECT 55.800 96.200 56.100 101.800 ;
        RECT 56.600 97.800 57.000 98.200 ;
        RECT 54.200 95.800 54.600 96.200 ;
        RECT 55.800 95.800 56.200 96.200 ;
        RECT 53.400 93.800 53.800 94.200 ;
        RECT 55.800 93.800 56.200 94.200 ;
        RECT 49.400 93.100 49.800 93.500 ;
        RECT 50.100 93.200 52.200 93.500 ;
        RECT 52.700 93.100 53.100 93.500 ;
        RECT 55.800 92.200 56.100 93.800 ;
        RECT 48.600 91.800 49.000 92.200 ;
        RECT 54.200 91.800 54.600 92.200 ;
        RECT 55.800 91.800 56.200 92.200 ;
        RECT 48.600 87.200 48.900 91.800 ;
        RECT 51.800 89.800 52.200 90.200 ;
        RECT 51.800 89.200 52.100 89.800 ;
        RECT 51.800 88.800 52.200 89.200 ;
        RECT 49.500 87.800 49.900 87.900 ;
        RECT 49.500 87.500 52.300 87.800 ;
        RECT 52.600 87.500 53.000 87.900 ;
        RECT 47.800 86.800 48.200 87.200 ;
        RECT 48.600 86.800 49.000 87.200 ;
        RECT 42.200 86.100 42.600 86.200 ;
        RECT 43.000 86.100 43.400 86.200 ;
        RECT 42.200 85.800 43.400 86.100 ;
        RECT 46.200 85.800 46.600 86.200 ;
        RECT 47.000 85.800 47.400 86.200 ;
        RECT 46.200 85.200 46.500 85.800 ;
        RECT 40.600 84.800 41.000 85.200 ;
        RECT 41.400 84.800 41.800 85.200 ;
        RECT 43.000 84.800 43.400 85.200 ;
        RECT 46.200 84.800 46.600 85.200 ;
        RECT 41.400 84.200 41.700 84.800 ;
        RECT 43.000 84.200 43.300 84.800 ;
        RECT 41.400 83.800 41.800 84.200 ;
        RECT 43.000 83.800 43.400 84.200 ;
        RECT 42.200 80.800 42.600 81.200 ;
        RECT 42.200 79.200 42.500 80.800 ;
        RECT 39.000 78.800 39.400 79.200 ;
        RECT 42.200 78.800 42.600 79.200 ;
        RECT 37.400 75.000 37.800 75.100 ;
        RECT 38.200 75.000 38.600 75.100 ;
        RECT 37.400 74.700 38.600 75.000 ;
        RECT 36.600 73.800 37.000 74.200 ;
        RECT 37.400 73.800 37.800 74.200 ;
        RECT 33.400 68.800 33.800 69.200 ;
        RECT 37.400 67.200 37.700 73.800 ;
        RECT 39.000 72.100 39.400 77.900 ;
        RECT 45.400 76.800 45.800 77.200 ;
        RECT 45.400 76.200 45.700 76.800 ;
        RECT 39.800 72.800 40.200 73.200 ;
        RECT 40.600 73.100 41.000 75.900 ;
        RECT 43.000 75.800 43.400 76.200 ;
        RECT 45.400 75.800 45.800 76.200 ;
        RECT 43.000 75.200 43.300 75.800 ;
        RECT 47.800 75.200 48.100 86.800 ;
        RECT 49.500 85.100 49.800 87.500 ;
        RECT 50.200 87.400 50.600 87.500 ;
        RECT 51.900 87.400 52.300 87.500 ;
        RECT 52.700 87.100 53.000 87.500 ;
        RECT 50.200 86.800 53.000 87.100 ;
        RECT 53.400 87.800 53.800 88.200 ;
        RECT 53.400 87.200 53.700 87.800 ;
        RECT 53.400 86.800 53.800 87.200 ;
        RECT 50.200 86.100 50.500 86.800 ;
        RECT 50.100 85.700 50.500 86.100 ;
        RECT 52.700 85.100 53.000 86.800 ;
        RECT 49.500 84.700 49.900 85.100 ;
        RECT 52.600 84.700 53.000 85.100 ;
        RECT 54.200 85.200 54.500 91.800 ;
        RECT 56.600 86.200 56.900 97.800 ;
        RECT 58.200 95.200 58.500 113.800 ;
        RECT 60.600 113.200 60.900 114.800 ;
        RECT 61.400 114.200 61.700 114.800 ;
        RECT 61.400 113.800 61.800 114.200 ;
        RECT 63.000 113.800 63.400 114.200 ;
        RECT 63.000 113.200 63.300 113.800 ;
        RECT 60.600 112.800 61.000 113.200 ;
        RECT 63.000 113.100 63.400 113.200 ;
        RECT 63.800 113.100 64.100 126.800 ;
        RECT 65.400 124.200 65.700 127.800 ;
        RECT 67.800 127.100 68.200 127.200 ;
        RECT 66.200 126.800 68.200 127.100 ;
        RECT 66.200 126.200 66.500 126.800 ;
        RECT 69.400 126.200 69.700 133.800 ;
        RECT 71.000 133.200 71.300 133.800 ;
        RECT 75.000 133.200 75.300 133.800 ;
        RECT 75.700 133.500 76.000 135.900 ;
        RECT 77.000 134.200 77.400 134.300 ;
        RECT 79.100 134.200 79.400 135.900 ;
        RECT 80.600 135.200 80.900 143.800 ;
        RECT 81.400 143.100 81.800 148.900 ;
        RECT 87.800 148.800 88.200 149.200 ;
        RECT 82.200 147.800 82.600 148.200 ;
        RECT 83.800 148.100 84.200 148.200 ;
        RECT 84.600 148.100 85.000 148.200 ;
        RECT 82.200 147.200 82.500 147.800 ;
        RECT 82.200 146.800 82.600 147.200 ;
        RECT 83.000 145.100 83.400 147.900 ;
        RECT 83.800 147.800 85.000 148.100 ;
        RECT 88.600 147.200 88.900 153.800 ;
        RECT 89.400 153.100 89.800 155.900 ;
        RECT 90.200 153.200 90.500 167.800 ;
        RECT 93.400 163.100 93.800 168.900 ;
        RECT 97.400 166.800 97.800 167.200 ;
        RECT 97.400 166.300 97.700 166.800 ;
        RECT 94.200 165.800 94.600 166.200 ;
        RECT 97.400 165.900 97.800 166.300 ;
        RECT 94.200 163.200 94.500 165.800 ;
        RECT 94.200 162.800 94.600 163.200 ;
        RECT 98.200 163.100 98.600 168.900 ;
        RECT 99.800 165.100 100.200 167.900 ;
        RECT 102.200 167.800 102.600 168.200 ;
        RECT 100.600 166.100 101.000 166.200 ;
        RECT 101.400 166.100 101.800 166.200 ;
        RECT 100.600 165.800 101.800 166.100 ;
        RECT 102.200 165.200 102.500 167.800 ;
        RECT 103.800 165.800 104.200 166.200 ;
        RECT 103.800 165.200 104.100 165.800 ;
        RECT 102.200 164.800 102.600 165.200 ;
        RECT 103.800 164.800 104.200 165.200 ;
        RECT 109.400 163.100 109.800 168.900 ;
        RECT 111.800 166.100 112.200 166.200 ;
        RECT 112.600 166.100 113.000 166.200 ;
        RECT 111.800 165.800 113.000 166.100 ;
        RECT 111.800 164.800 112.200 165.200 ;
        RECT 91.000 162.100 91.400 162.200 ;
        RECT 91.800 162.100 92.200 162.200 ;
        RECT 91.000 161.800 92.200 162.100 ;
        RECT 107.000 162.100 107.400 162.200 ;
        RECT 107.800 162.100 108.200 162.200 ;
        RECT 107.000 161.800 108.200 162.100 ;
        RECT 111.000 161.800 111.400 162.200 ;
        RECT 98.200 157.100 98.600 157.200 ;
        RECT 99.000 157.100 99.400 157.200 ;
        RECT 98.200 156.800 99.400 157.100 ;
        RECT 103.000 156.800 103.400 157.200 ;
        RECT 91.000 155.800 91.400 156.200 ;
        RECT 95.000 155.800 95.400 156.200 ;
        RECT 101.400 156.100 101.800 156.200 ;
        RECT 102.200 156.100 102.600 156.200 ;
        RECT 101.400 155.800 102.600 156.100 ;
        RECT 91.000 155.200 91.300 155.800 ;
        RECT 95.000 155.200 95.300 155.800 ;
        RECT 103.000 155.200 103.300 156.800 ;
        RECT 111.000 155.200 111.300 161.800 ;
        RECT 111.800 159.200 112.100 164.800 ;
        RECT 114.200 163.100 114.600 168.900 ;
        RECT 115.000 167.800 115.400 168.200 ;
        RECT 115.000 167.200 115.300 167.800 ;
        RECT 115.000 166.800 115.400 167.200 ;
        RECT 115.800 165.100 116.200 167.900 ;
        RECT 118.200 165.800 118.600 166.200 ;
        RECT 119.000 165.800 119.400 166.200 ;
        RECT 111.800 158.800 112.200 159.200 ;
        RECT 118.200 156.200 118.500 165.800 ;
        RECT 119.000 160.200 119.300 165.800 ;
        RECT 123.800 163.100 124.200 168.900 ;
        RECT 127.000 166.800 127.400 167.200 ;
        RECT 127.000 166.200 127.300 166.800 ;
        RECT 124.600 165.800 125.000 166.200 ;
        RECT 127.000 165.800 127.400 166.200 ;
        RECT 124.600 163.200 124.900 165.800 ;
        RECT 124.600 162.800 125.000 163.200 ;
        RECT 128.600 163.100 129.000 168.900 ;
        RECT 130.200 165.100 130.600 167.900 ;
        RECT 135.800 165.100 136.200 167.900 ;
        RECT 137.400 163.100 137.800 168.900 ;
        RECT 138.200 167.800 138.600 168.200 ;
        RECT 138.200 167.200 138.500 167.800 ;
        RECT 138.200 166.800 138.600 167.200 ;
        RECT 139.000 166.800 139.400 167.200 ;
        RECT 121.400 161.800 121.800 162.200 ;
        RECT 119.000 159.800 119.400 160.200 ;
        RECT 121.400 158.200 121.700 161.800 ;
        RECT 127.000 159.800 127.400 160.200 ;
        RECT 129.400 159.800 129.800 160.200 ;
        RECT 127.000 159.200 127.300 159.800 ;
        RECT 127.000 158.800 127.400 159.200 ;
        RECT 121.400 157.800 121.800 158.200 ;
        RECT 118.200 155.800 118.600 156.200 ;
        RECT 123.800 155.800 124.200 156.200 ;
        RECT 128.600 155.800 129.000 156.200 ;
        RECT 123.800 155.200 124.100 155.800 ;
        RECT 128.600 155.200 128.900 155.800 ;
        RECT 129.400 155.200 129.700 159.800 ;
        RECT 131.000 157.800 131.400 158.200 ;
        RECT 91.000 154.800 91.400 155.200 ;
        RECT 94.200 154.800 94.600 155.200 ;
        RECT 95.000 154.800 95.400 155.200 ;
        RECT 95.800 154.800 96.200 155.200 ;
        RECT 99.800 155.100 100.200 155.200 ;
        RECT 100.600 155.100 101.000 155.200 ;
        RECT 99.800 154.800 101.000 155.100 ;
        RECT 101.400 155.100 101.800 155.200 ;
        RECT 102.200 155.100 102.600 155.200 ;
        RECT 101.400 154.800 102.600 155.100 ;
        RECT 103.000 154.800 103.400 155.200 ;
        RECT 107.800 155.100 108.200 155.200 ;
        RECT 108.600 155.100 109.000 155.200 ;
        RECT 107.800 154.800 109.000 155.100 ;
        RECT 110.200 154.800 110.600 155.200 ;
        RECT 111.000 154.800 111.400 155.200 ;
        RECT 113.400 154.800 113.800 155.200 ;
        RECT 115.000 154.800 115.400 155.200 ;
        RECT 121.400 155.100 121.800 155.200 ;
        RECT 122.200 155.100 122.600 155.200 ;
        RECT 121.400 154.800 122.600 155.100 ;
        RECT 123.800 154.800 124.200 155.200 ;
        RECT 125.400 155.100 125.800 155.200 ;
        RECT 126.200 155.100 126.600 155.200 ;
        RECT 125.400 154.800 126.600 155.100 ;
        RECT 127.800 154.800 128.200 155.200 ;
        RECT 128.600 154.800 129.000 155.200 ;
        RECT 129.400 154.800 129.800 155.200 ;
        RECT 130.200 154.800 130.600 155.200 ;
        RECT 92.600 153.800 93.000 154.200 ;
        RECT 92.600 153.200 92.900 153.800 ;
        RECT 90.200 152.800 90.600 153.200 ;
        RECT 92.600 152.800 93.000 153.200 ;
        RECT 91.000 148.800 91.400 149.200 ;
        RECT 83.800 146.800 84.200 147.200 ;
        RECT 86.200 147.100 86.600 147.200 ;
        RECT 87.000 147.100 87.400 147.200 ;
        RECT 86.200 146.800 87.400 147.100 ;
        RECT 88.600 146.800 89.000 147.200 ;
        RECT 83.800 146.200 84.100 146.800 ;
        RECT 91.000 146.200 91.300 148.800 ;
        RECT 91.800 146.800 92.200 147.200 ;
        RECT 91.800 146.200 92.100 146.800 ;
        RECT 94.200 146.200 94.500 154.800 ;
        RECT 95.000 149.200 95.300 154.800 ;
        RECT 95.800 154.200 96.100 154.800 ;
        RECT 95.800 153.800 96.200 154.200 ;
        RECT 96.600 153.100 97.000 153.200 ;
        RECT 97.400 153.100 97.800 153.200 ;
        RECT 96.600 152.800 97.800 153.100 ;
        RECT 101.400 152.800 101.800 153.200 ;
        RECT 103.800 153.100 104.200 153.200 ;
        RECT 104.600 153.100 105.000 153.200 ;
        RECT 103.800 152.800 105.000 153.100 ;
        RECT 108.600 152.800 109.000 153.200 ;
        RECT 101.400 149.200 101.700 152.800 ;
        RECT 95.000 148.800 95.400 149.200 ;
        RECT 101.400 148.800 101.800 149.200 ;
        RECT 103.800 149.100 104.200 149.200 ;
        RECT 104.600 149.100 105.000 149.200 ;
        RECT 103.800 148.800 105.000 149.100 ;
        RECT 103.000 147.800 103.400 148.200 ;
        RECT 103.800 147.800 104.200 148.200 ;
        RECT 83.800 145.800 84.200 146.200 ;
        RECT 85.400 145.800 85.800 146.200 ;
        RECT 86.200 146.100 86.600 146.200 ;
        RECT 87.000 146.100 87.400 146.200 ;
        RECT 86.200 145.800 87.400 146.100 ;
        RECT 91.000 145.800 91.400 146.200 ;
        RECT 91.800 145.800 92.200 146.200 ;
        RECT 93.400 145.800 93.800 146.200 ;
        RECT 94.200 145.800 94.600 146.200 ;
        RECT 96.600 145.800 97.000 146.200 ;
        RECT 99.000 145.800 99.400 146.200 ;
        RECT 85.400 144.200 85.700 145.800 ;
        RECT 83.000 143.800 83.400 144.200 ;
        RECT 85.400 143.800 85.800 144.200 ;
        RECT 81.400 141.800 81.800 142.200 ;
        RECT 81.400 135.200 81.700 141.800 ;
        RECT 83.000 139.200 83.300 143.800 ;
        RECT 86.200 143.200 86.500 145.800 ;
        RECT 88.600 145.100 89.000 145.200 ;
        RECT 89.400 145.100 89.800 145.200 ;
        RECT 88.600 144.800 89.800 145.100 ;
        RECT 86.200 142.800 86.600 143.200 ;
        RECT 83.000 138.800 83.400 139.200 ;
        RECT 88.600 136.200 88.900 144.800 ;
        RECT 90.200 142.800 90.600 143.200 ;
        RECT 90.200 141.200 90.500 142.800 ;
        RECT 90.200 140.800 90.600 141.200 ;
        RECT 88.600 135.800 89.000 136.200 ;
        RECT 80.600 134.800 81.000 135.200 ;
        RECT 81.400 134.800 81.800 135.200 ;
        RECT 83.800 134.800 84.200 135.200 ;
        RECT 84.600 134.800 85.000 135.200 ;
        RECT 85.400 134.800 85.800 135.200 ;
        RECT 77.000 133.900 79.400 134.200 ;
        RECT 76.600 133.500 77.000 133.600 ;
        RECT 78.300 133.500 78.700 133.600 ;
        RECT 79.100 133.500 79.400 133.900 ;
        RECT 71.000 132.800 71.400 133.200 ;
        RECT 75.000 132.800 75.400 133.200 ;
        RECT 75.700 133.100 76.100 133.500 ;
        RECT 76.600 133.200 78.700 133.500 ;
        RECT 66.200 125.800 66.600 126.200 ;
        RECT 67.000 125.800 67.400 126.200 ;
        RECT 67.800 125.800 68.200 126.200 ;
        RECT 69.400 125.800 69.800 126.200 ;
        RECT 67.000 125.200 67.300 125.800 ;
        RECT 67.800 125.200 68.100 125.800 ;
        RECT 67.000 124.800 67.400 125.200 ;
        RECT 67.800 124.800 68.200 125.200 ;
        RECT 65.400 123.800 65.800 124.200 ;
        RECT 67.000 123.200 67.300 124.800 ;
        RECT 67.000 122.800 67.400 123.200 ;
        RECT 69.400 122.800 69.800 123.200 ;
        RECT 69.400 119.200 69.700 122.800 ;
        RECT 69.400 118.800 69.800 119.200 ;
        RECT 65.400 116.800 65.800 117.200 ;
        RECT 68.600 116.800 69.000 117.200 ;
        RECT 65.400 115.200 65.700 116.800 ;
        RECT 68.600 115.200 68.900 116.800 ;
        RECT 71.000 115.200 71.300 132.800 ;
        RECT 71.800 131.800 72.200 132.200 ;
        RECT 71.800 129.200 72.100 131.800 ;
        RECT 71.800 128.800 72.200 129.200 ;
        RECT 72.600 128.800 73.000 129.200 ;
        RECT 72.600 128.200 72.900 128.800 ;
        RECT 71.800 127.800 72.200 128.200 ;
        RECT 72.600 127.800 73.000 128.200 ;
        RECT 76.600 127.800 77.000 128.200 ;
        RECT 71.800 127.200 72.100 127.800 ;
        RECT 71.800 126.800 72.200 127.200 ;
        RECT 72.600 125.800 73.000 126.200 ;
        RECT 72.600 125.200 72.900 125.800 ;
        RECT 72.600 124.800 73.000 125.200 ;
        RECT 76.600 123.200 76.900 127.800 ;
        RECT 78.200 127.200 78.500 133.200 ;
        RECT 79.000 133.100 79.400 133.500 ;
        RECT 79.800 133.800 80.200 134.200 ;
        RECT 79.800 127.200 80.100 133.800 ;
        RECT 78.200 126.800 78.600 127.200 ;
        RECT 79.800 126.800 80.200 127.200 ;
        RECT 79.800 126.200 80.100 126.800 ;
        RECT 79.800 125.800 80.200 126.200 ;
        RECT 79.800 124.800 80.200 125.200 ;
        RECT 79.800 124.200 80.100 124.800 ;
        RECT 77.400 124.100 77.800 124.200 ;
        RECT 78.200 124.100 78.600 124.200 ;
        RECT 77.400 123.800 78.600 124.100 ;
        RECT 79.800 123.800 80.200 124.200 ;
        RECT 76.600 122.800 77.000 123.200 ;
        RECT 65.400 114.800 65.800 115.200 ;
        RECT 68.600 114.800 69.000 115.200 ;
        RECT 71.000 114.800 71.400 115.200 ;
        RECT 63.000 112.800 64.100 113.100 ;
        RECT 67.000 112.800 67.400 113.200 ;
        RECT 68.600 112.800 69.000 113.200 ;
        RECT 62.200 110.800 62.600 111.200 ;
        RECT 61.400 107.800 61.800 108.200 ;
        RECT 61.400 107.200 61.700 107.800 ;
        RECT 59.000 106.800 59.400 107.200 ;
        RECT 61.400 106.800 61.800 107.200 ;
        RECT 59.000 106.200 59.300 106.800 ;
        RECT 62.200 106.200 62.500 110.800 ;
        RECT 59.000 105.800 59.400 106.200 ;
        RECT 62.200 105.800 62.600 106.200 ;
        RECT 59.000 105.100 59.400 105.200 ;
        RECT 59.800 105.100 60.200 105.200 ;
        RECT 59.000 104.800 60.200 105.100 ;
        RECT 60.600 104.800 61.000 105.200 ;
        RECT 60.600 104.200 60.900 104.800 ;
        RECT 60.600 103.800 61.000 104.200 ;
        RECT 60.600 98.200 60.900 103.800 ;
        RECT 62.200 101.800 62.600 102.200 ;
        RECT 60.600 97.800 61.000 98.200 ;
        RECT 62.200 95.200 62.500 101.800 ;
        RECT 58.200 94.800 58.600 95.200 ;
        RECT 59.000 95.100 59.400 95.200 ;
        RECT 59.800 95.100 60.200 95.200 ;
        RECT 59.000 94.800 60.200 95.100 ;
        RECT 61.400 94.800 61.800 95.200 ;
        RECT 62.200 94.800 62.600 95.200 ;
        RECT 57.400 93.800 57.800 94.200 ;
        RECT 57.400 90.200 57.700 93.800 ;
        RECT 61.400 93.200 61.700 94.800 ;
        RECT 63.000 94.200 63.300 112.800 ;
        RECT 67.000 112.200 67.300 112.800 ;
        RECT 63.800 111.800 64.200 112.200 ;
        RECT 66.200 111.800 66.600 112.200 ;
        RECT 67.000 111.800 67.400 112.200 ;
        RECT 67.800 111.800 68.200 112.200 ;
        RECT 63.800 108.200 64.100 111.800 ;
        RECT 66.200 109.200 66.500 111.800 ;
        RECT 67.800 111.200 68.100 111.800 ;
        RECT 67.800 110.800 68.200 111.200 ;
        RECT 66.200 108.800 66.600 109.200 ;
        RECT 63.800 107.800 64.200 108.200 ;
        RECT 64.600 107.800 65.000 108.200 ;
        RECT 65.400 107.800 65.800 108.200 ;
        RECT 64.600 107.200 64.900 107.800 ;
        RECT 65.400 107.200 65.700 107.800 ;
        RECT 64.600 106.800 65.000 107.200 ;
        RECT 65.400 106.800 65.800 107.200 ;
        RECT 67.000 107.100 67.400 107.200 ;
        RECT 67.800 107.100 68.200 107.200 ;
        RECT 67.000 106.800 68.200 107.100 ;
        RECT 68.600 107.000 68.900 112.800 ;
        RECT 71.800 112.100 72.200 117.900 ;
        RECT 75.800 117.800 76.200 118.200 ;
        RECT 75.800 115.100 76.100 117.800 ;
        RECT 75.800 114.700 76.200 115.100 ;
        RECT 76.600 112.100 77.000 117.900 ;
        RECT 79.800 116.800 80.200 117.200 ;
        RECT 77.400 113.800 77.800 114.200 ;
        RECT 77.400 113.200 77.700 113.800 ;
        RECT 77.400 112.800 77.800 113.200 ;
        RECT 78.200 113.100 78.600 115.900 ;
        RECT 79.800 113.200 80.100 116.800 ;
        RECT 80.600 116.200 80.900 134.800 ;
        RECT 81.400 120.200 81.700 134.800 ;
        RECT 83.800 132.200 84.100 134.800 ;
        RECT 84.600 134.200 84.900 134.800 ;
        RECT 85.400 134.200 85.700 134.800 ;
        RECT 84.600 133.800 85.000 134.200 ;
        RECT 85.400 133.800 85.800 134.200 ;
        RECT 83.800 131.800 84.200 132.200 ;
        RECT 87.000 131.800 87.400 132.200 ;
        RECT 83.800 130.200 84.100 131.800 ;
        RECT 83.800 129.800 84.200 130.200 ;
        RECT 82.200 129.100 82.600 129.200 ;
        RECT 83.000 129.100 83.400 129.200 ;
        RECT 82.200 128.800 83.400 129.100 ;
        RECT 83.800 127.800 84.200 128.200 ;
        RECT 83.800 127.200 84.100 127.800 ;
        RECT 83.800 126.800 84.200 127.200 ;
        RECT 82.200 125.100 82.600 125.200 ;
        RECT 83.000 125.100 83.400 125.200 ;
        RECT 82.200 124.800 83.400 125.100 ;
        RECT 81.400 119.800 81.800 120.200 ;
        RECT 83.800 117.200 84.100 126.800 ;
        RECT 87.000 126.200 87.300 131.800 ;
        RECT 88.600 131.200 88.900 135.800 ;
        RECT 90.200 135.200 90.500 140.800 ;
        RECT 90.200 134.800 90.600 135.200 ;
        RECT 87.800 130.800 88.200 131.200 ;
        RECT 88.600 130.800 89.000 131.200 ;
        RECT 87.800 129.200 88.100 130.800 ;
        RECT 87.800 128.800 88.200 129.200 ;
        RECT 84.600 126.100 85.000 126.200 ;
        RECT 85.400 126.100 85.800 126.200 ;
        RECT 84.600 125.800 85.800 126.100 ;
        RECT 87.000 125.800 87.400 126.200 ;
        RECT 88.600 125.800 89.000 126.200 ;
        RECT 87.000 118.200 87.300 125.800 ;
        RECT 88.600 125.200 88.900 125.800 ;
        RECT 88.600 124.800 89.000 125.200 ;
        RECT 87.000 117.800 87.400 118.200 ;
        RECT 83.800 116.800 84.200 117.200 ;
        RECT 80.600 115.800 81.000 116.200 ;
        RECT 83.800 115.800 84.200 116.200 ;
        RECT 86.200 115.800 86.600 116.200 ;
        RECT 83.800 115.200 84.100 115.800 ;
        RECT 86.200 115.200 86.500 115.800 ;
        RECT 81.400 114.800 81.800 115.200 ;
        RECT 83.800 114.800 84.200 115.200 ;
        RECT 86.200 114.800 86.600 115.200 ;
        RECT 87.000 114.800 87.400 115.200 ;
        RECT 89.400 114.800 89.800 115.200 ;
        RECT 81.400 114.200 81.700 114.800 ;
        RECT 81.400 113.800 81.800 114.200 ;
        RECT 79.800 112.800 80.200 113.200 ;
        RECT 76.600 109.800 77.000 110.200 ;
        RECT 76.600 109.200 76.900 109.800 ;
        RECT 70.200 108.800 70.600 109.200 ;
        RECT 76.600 108.800 77.000 109.200 ;
        RECT 82.200 109.100 82.600 109.200 ;
        RECT 83.000 109.100 83.400 109.200 ;
        RECT 82.200 108.800 83.400 109.100 ;
        RECT 83.800 109.100 84.100 114.800 ;
        RECT 85.400 114.100 85.800 114.200 ;
        RECT 86.200 114.100 86.600 114.200 ;
        RECT 85.400 113.800 86.600 114.100 ;
        RECT 85.400 112.200 85.700 113.800 ;
        RECT 85.400 111.800 85.800 112.200 ;
        RECT 87.000 110.200 87.300 114.800 ;
        RECT 89.400 111.200 89.700 114.800 ;
        RECT 89.400 110.800 89.800 111.200 ;
        RECT 90.200 110.200 90.500 134.800 ;
        RECT 91.800 134.200 92.100 145.800 ;
        RECT 93.400 143.200 93.700 145.800 ;
        RECT 94.200 144.800 94.600 145.200 ;
        RECT 93.400 142.800 93.800 143.200 ;
        RECT 94.200 139.200 94.500 144.800 ;
        RECT 94.200 138.800 94.600 139.200 ;
        RECT 96.600 135.200 96.900 145.800 ;
        RECT 92.600 135.100 93.000 135.200 ;
        RECT 93.400 135.100 93.800 135.200 ;
        RECT 92.600 134.800 93.800 135.100 ;
        RECT 96.600 134.800 97.000 135.200 ;
        RECT 91.000 134.100 91.400 134.200 ;
        RECT 91.800 134.100 92.200 134.200 ;
        RECT 91.000 133.800 92.200 134.100 ;
        RECT 91.000 123.800 91.400 124.200 ;
        RECT 91.000 123.200 91.300 123.800 ;
        RECT 91.000 122.800 91.400 123.200 ;
        RECT 93.400 123.100 93.800 128.900 ;
        RECT 95.800 126.100 96.200 126.200 ;
        RECT 96.600 126.100 97.000 126.200 ;
        RECT 95.800 125.800 97.000 126.100 ;
        RECT 98.200 123.100 98.600 128.900 ;
        RECT 99.000 127.200 99.300 145.800 ;
        RECT 100.600 137.800 101.000 138.200 ;
        RECT 100.600 135.200 100.900 137.800 ;
        RECT 101.400 135.800 101.800 136.200 ;
        RECT 101.400 135.200 101.700 135.800 ;
        RECT 100.600 134.800 101.000 135.200 ;
        RECT 101.400 134.800 101.800 135.200 ;
        RECT 99.000 126.800 99.400 127.200 ;
        RECT 91.000 112.800 91.400 113.200 ;
        RECT 92.600 113.100 93.000 113.200 ;
        RECT 93.400 113.100 93.800 113.200 ;
        RECT 92.600 112.800 93.800 113.100 ;
        RECT 87.000 109.800 87.400 110.200 ;
        RECT 90.200 109.800 90.600 110.200 ;
        RECT 87.000 109.200 87.300 109.800 ;
        RECT 83.800 108.800 84.900 109.100 ;
        RECT 70.200 108.200 70.500 108.800 ;
        RECT 70.200 107.800 70.600 108.200 ;
        RECT 75.000 107.800 75.400 108.200 ;
        RECT 77.400 107.800 77.800 108.200 ;
        RECT 68.600 106.600 69.000 107.000 ;
        RECT 68.600 106.200 68.900 106.600 ;
        RECT 75.000 106.200 75.300 107.800 ;
        RECT 63.800 106.100 64.200 106.200 ;
        RECT 64.600 106.100 65.000 106.200 ;
        RECT 63.800 105.800 65.000 106.100 ;
        RECT 65.400 106.100 65.800 106.200 ;
        RECT 66.200 106.100 66.600 106.200 ;
        RECT 65.400 105.800 66.600 106.100 ;
        RECT 67.000 106.100 67.400 106.200 ;
        RECT 67.800 106.100 68.200 106.200 ;
        RECT 67.000 105.800 68.200 106.100 ;
        RECT 68.600 105.800 69.000 106.200 ;
        RECT 73.400 105.800 73.800 106.200 ;
        RECT 75.000 105.800 75.400 106.200 ;
        RECT 70.200 105.100 70.600 105.200 ;
        RECT 71.000 105.100 71.400 105.200 ;
        RECT 70.200 104.800 71.400 105.100 ;
        RECT 73.400 104.200 73.700 105.800 ;
        RECT 73.400 103.800 73.800 104.200 ;
        RECT 77.400 103.200 77.700 107.800 ;
        RECT 83.800 105.800 84.200 106.200 ;
        RECT 77.400 102.800 77.800 103.200 ;
        RECT 73.400 100.800 73.800 101.200 ;
        RECT 63.800 95.900 64.200 96.300 ;
        RECT 66.900 95.900 67.300 96.300 ;
        RECT 73.400 96.200 73.700 100.800 ;
        RECT 63.800 94.200 64.100 95.900 ;
        RECT 66.300 94.900 66.700 95.300 ;
        RECT 66.300 94.200 66.600 94.900 ;
        RECT 63.000 93.800 63.400 94.200 ;
        RECT 63.800 93.900 66.600 94.200 ;
        RECT 63.000 93.200 63.300 93.800 ;
        RECT 63.800 93.500 64.100 93.900 ;
        RECT 64.500 93.500 64.900 93.600 ;
        RECT 66.200 93.500 66.600 93.600 ;
        RECT 67.000 93.500 67.300 95.900 ;
        RECT 72.600 95.800 73.000 96.200 ;
        RECT 73.400 95.800 73.800 96.200 ;
        RECT 58.200 93.100 58.600 93.200 ;
        RECT 59.000 93.100 59.400 93.200 ;
        RECT 58.200 92.800 59.400 93.100 ;
        RECT 61.400 92.800 61.800 93.200 ;
        RECT 63.000 92.800 63.400 93.200 ;
        RECT 63.800 93.100 64.200 93.500 ;
        RECT 64.500 93.200 67.300 93.500 ;
        RECT 66.900 93.100 67.300 93.200 ;
        RECT 67.800 94.800 68.200 95.200 ;
        RECT 71.000 94.800 71.400 95.200 ;
        RECT 67.800 94.200 68.100 94.800 ;
        RECT 67.800 93.800 68.200 94.200 ;
        RECT 68.600 93.800 69.000 94.200 ;
        RECT 58.200 91.800 58.600 92.200 ;
        RECT 58.200 91.200 58.500 91.800 ;
        RECT 58.200 90.800 58.600 91.200 ;
        RECT 57.400 89.800 57.800 90.200 ;
        RECT 67.800 89.200 68.100 93.800 ;
        RECT 68.600 93.200 68.900 93.800 ;
        RECT 68.600 92.800 69.000 93.200 ;
        RECT 71.000 93.100 71.300 94.800 ;
        RECT 71.000 92.800 72.100 93.100 ;
        RECT 58.200 88.800 58.600 89.200 ;
        RECT 62.200 89.100 62.600 89.200 ;
        RECT 63.000 89.100 63.400 89.200 ;
        RECT 62.200 88.800 63.400 89.100 ;
        RECT 58.200 88.200 58.500 88.800 ;
        RECT 58.200 87.800 58.600 88.200 ;
        RECT 56.600 85.800 57.000 86.200 ;
        RECT 59.800 86.100 60.200 86.200 ;
        RECT 60.600 86.100 61.000 86.200 ;
        RECT 59.800 85.800 61.000 86.100 ;
        RECT 54.200 84.800 54.600 85.200 ;
        RECT 59.000 84.800 59.400 85.200 ;
        RECT 59.000 84.200 59.300 84.800 ;
        RECT 59.000 83.800 59.400 84.200 ;
        RECT 59.800 83.800 60.200 84.200 ;
        RECT 59.800 79.200 60.100 83.800 ;
        RECT 64.600 83.100 65.000 88.900 ;
        RECT 67.800 88.800 68.200 89.200 ;
        RECT 68.600 86.800 69.000 87.200 ;
        RECT 68.600 86.300 68.900 86.800 ;
        RECT 66.200 85.800 66.600 86.200 ;
        RECT 68.600 85.900 69.000 86.300 ;
        RECT 61.400 81.800 61.800 82.200 ;
        RECT 59.800 78.800 60.200 79.200 ;
        RECT 48.600 76.800 49.000 77.200 ;
        RECT 51.000 76.800 51.400 77.200 ;
        RECT 55.800 76.800 56.200 77.200 ;
        RECT 42.200 74.800 42.600 75.200 ;
        RECT 43.000 74.800 43.400 75.200 ;
        RECT 47.800 74.800 48.200 75.200 ;
        RECT 41.400 72.800 41.800 73.200 ;
        RECT 38.200 69.800 38.600 70.200 ;
        RECT 38.200 68.200 38.500 69.800 ;
        RECT 38.200 67.800 38.600 68.200 ;
        RECT 37.400 66.800 37.800 67.200 ;
        RECT 36.600 65.800 37.000 66.200 ;
        RECT 33.400 65.100 33.800 65.200 ;
        RECT 34.200 65.100 34.600 65.200 ;
        RECT 33.400 64.800 34.600 65.100 ;
        RECT 36.600 62.200 36.900 65.800 ;
        RECT 36.600 62.100 37.000 62.200 ;
        RECT 36.600 61.800 37.700 62.100 ;
        RECT 35.000 59.800 35.400 60.200 ;
        RECT 27.800 54.800 28.200 55.200 ;
        RECT 27.800 53.800 28.200 54.200 ;
        RECT 30.200 53.800 30.600 54.200 ;
        RECT 27.800 53.200 28.100 53.800 ;
        RECT 30.200 53.200 30.500 53.800 ;
        RECT 31.100 53.500 31.400 55.900 ;
        RECT 31.800 55.800 32.200 56.200 ;
        RECT 34.200 55.900 34.600 56.300 ;
        RECT 31.700 54.900 32.100 55.300 ;
        RECT 31.800 54.200 32.100 54.900 ;
        RECT 34.300 54.200 34.600 55.900 ;
        RECT 31.800 53.900 34.600 54.200 ;
        RECT 31.800 53.500 32.200 53.600 ;
        RECT 33.500 53.500 33.900 53.600 ;
        RECT 34.300 53.500 34.600 53.900 ;
        RECT 35.000 54.200 35.300 59.800 ;
        RECT 37.400 56.200 37.700 61.800 ;
        RECT 38.200 60.200 38.500 67.800 ;
        RECT 39.000 65.100 39.400 67.900 ;
        RECT 39.800 67.200 40.100 72.800 ;
        RECT 39.800 66.800 40.200 67.200 ;
        RECT 40.600 63.100 41.000 68.900 ;
        RECT 41.400 66.200 41.700 72.800 ;
        RECT 42.200 71.200 42.500 74.800 ;
        RECT 43.000 74.100 43.400 74.200 ;
        RECT 43.800 74.100 44.200 74.200 ;
        RECT 43.000 73.800 44.200 74.100 ;
        RECT 47.000 73.100 47.400 73.200 ;
        RECT 47.800 73.100 48.200 73.200 ;
        RECT 47.000 72.800 48.200 73.100 ;
        RECT 42.200 70.800 42.600 71.200 ;
        RECT 42.200 66.200 42.500 70.800 ;
        RECT 48.600 69.200 48.900 76.800 ;
        RECT 51.000 76.200 51.300 76.800 ;
        RECT 55.800 76.200 56.100 76.800 ;
        RECT 51.000 75.800 51.400 76.200 ;
        RECT 51.800 75.800 52.200 76.200 ;
        RECT 53.400 76.100 53.800 76.200 ;
        RECT 54.200 76.100 54.600 76.200 ;
        RECT 53.400 75.800 54.600 76.100 ;
        RECT 55.800 75.800 56.200 76.200 ;
        RECT 49.400 75.100 49.800 75.200 ;
        RECT 51.800 75.100 52.100 75.800 ;
        RECT 49.400 74.800 52.100 75.100 ;
        RECT 55.800 74.800 56.200 75.200 ;
        RECT 56.600 74.800 57.000 75.200 ;
        RECT 59.800 75.100 60.200 75.200 ;
        RECT 60.600 75.100 61.000 75.200 ;
        RECT 59.800 74.800 61.000 75.100 ;
        RECT 55.800 74.200 56.100 74.800 ;
        RECT 56.600 74.200 56.900 74.800 ;
        RECT 53.400 73.800 53.800 74.200 ;
        RECT 55.800 73.800 56.200 74.200 ;
        RECT 56.600 73.800 57.000 74.200 ;
        RECT 57.400 74.100 57.800 74.200 ;
        RECT 58.200 74.100 58.600 74.200 ;
        RECT 57.400 73.800 58.600 74.100 ;
        RECT 53.400 73.200 53.700 73.800 ;
        RECT 59.800 73.200 60.100 74.800 ;
        RECT 61.400 74.200 61.700 81.800 ;
        RECT 65.400 77.800 65.800 78.200 ;
        RECT 65.400 77.200 65.700 77.800 ;
        RECT 64.600 77.100 65.000 77.200 ;
        RECT 63.800 76.800 65.000 77.100 ;
        RECT 65.400 76.800 65.800 77.200 ;
        RECT 61.400 73.800 61.800 74.200 ;
        RECT 63.000 73.800 63.400 74.200 ;
        RECT 63.000 73.200 63.300 73.800 ;
        RECT 49.400 73.100 49.800 73.200 ;
        RECT 50.200 73.100 50.600 73.200 ;
        RECT 49.400 72.800 50.600 73.100 ;
        RECT 51.000 73.100 51.400 73.200 ;
        RECT 51.800 73.100 52.200 73.200 ;
        RECT 51.000 72.800 52.200 73.100 ;
        RECT 53.400 72.800 53.800 73.200 ;
        RECT 57.400 72.800 57.800 73.200 ;
        RECT 59.800 72.800 60.200 73.200 ;
        RECT 63.000 72.800 63.400 73.200 ;
        RECT 52.600 71.800 53.000 72.200 ;
        RECT 41.400 65.800 41.800 66.200 ;
        RECT 42.200 65.800 42.600 66.200 ;
        RECT 43.000 65.800 43.400 66.200 ;
        RECT 38.200 59.800 38.600 60.200 ;
        RECT 35.800 55.800 36.200 56.200 ;
        RECT 37.400 55.800 37.800 56.200 ;
        RECT 39.800 56.100 40.200 56.200 ;
        RECT 40.600 56.100 41.000 56.200 ;
        RECT 39.800 55.800 41.000 56.100 ;
        RECT 35.000 53.800 35.400 54.200 ;
        RECT 31.100 53.200 33.900 53.500 ;
        RECT 27.800 52.800 28.200 53.200 ;
        RECT 30.200 52.800 30.600 53.200 ;
        RECT 31.100 53.100 31.500 53.200 ;
        RECT 34.200 53.100 34.600 53.500 ;
        RECT 35.800 53.200 36.100 55.800 ;
        RECT 37.400 55.200 37.700 55.800 ;
        RECT 37.400 54.800 37.800 55.200 ;
        RECT 42.200 53.800 42.600 54.200 ;
        RECT 42.200 53.200 42.500 53.800 ;
        RECT 43.000 53.200 43.300 65.800 ;
        RECT 45.400 63.100 45.800 68.900 ;
        RECT 48.600 68.800 49.000 69.200 ;
        RECT 52.600 68.200 52.900 71.800 ;
        RECT 53.400 70.200 53.700 72.800 ;
        RECT 53.400 69.800 53.800 70.200 ;
        RECT 50.200 67.800 50.600 68.200 ;
        RECT 52.600 67.800 53.000 68.200 ;
        RECT 50.200 66.200 50.500 67.800 ;
        RECT 53.400 67.200 53.700 69.800 ;
        RECT 55.000 67.800 55.400 68.200 ;
        RECT 55.000 67.200 55.300 67.800 ;
        RECT 53.400 66.800 53.800 67.200 ;
        RECT 54.200 66.800 54.600 67.200 ;
        RECT 55.000 66.800 55.400 67.200 ;
        RECT 56.600 66.800 57.000 67.200 ;
        RECT 54.200 66.200 54.500 66.800 ;
        RECT 56.600 66.200 56.900 66.800 ;
        RECT 50.200 65.800 50.600 66.200 ;
        RECT 53.400 65.800 53.800 66.200 ;
        RECT 54.200 65.800 54.600 66.200 ;
        RECT 56.600 65.800 57.000 66.200 ;
        RECT 53.400 65.200 53.700 65.800 ;
        RECT 57.400 65.200 57.700 72.800 ;
        RECT 59.800 71.800 60.200 72.200 ;
        RECT 62.200 71.800 62.600 72.200 ;
        RECT 59.800 67.200 60.100 71.800 ;
        RECT 62.200 71.200 62.500 71.800 ;
        RECT 62.200 70.800 62.600 71.200 ;
        RECT 63.000 69.800 63.400 70.200 ;
        RECT 63.000 69.200 63.300 69.800 ;
        RECT 62.200 68.800 62.600 69.200 ;
        RECT 63.000 68.800 63.400 69.200 ;
        RECT 62.200 68.200 62.500 68.800 ;
        RECT 63.800 68.200 64.100 76.800 ;
        RECT 66.200 76.200 66.500 85.800 ;
        RECT 69.400 83.100 69.800 88.900 ;
        RECT 70.200 86.800 70.600 87.200 ;
        RECT 65.400 75.800 65.800 76.200 ;
        RECT 66.200 75.800 66.600 76.200 ;
        RECT 65.400 75.200 65.700 75.800 ;
        RECT 65.400 74.800 65.800 75.200 ;
        RECT 64.600 71.800 65.000 72.200 ;
        RECT 67.000 71.800 67.400 72.200 ;
        RECT 69.400 72.100 69.800 77.900 ;
        RECT 70.200 75.200 70.500 86.800 ;
        RECT 71.000 85.100 71.400 87.900 ;
        RECT 71.800 85.200 72.100 92.800 ;
        RECT 72.600 89.200 72.900 95.800 ;
        RECT 73.400 95.200 73.700 95.800 ;
        RECT 77.400 95.200 77.700 102.800 ;
        RECT 81.400 97.800 81.800 98.200 ;
        RECT 80.600 95.800 81.000 96.200 ;
        RECT 80.600 95.200 80.900 95.800 ;
        RECT 81.400 95.200 81.700 97.800 ;
        RECT 83.800 95.200 84.100 105.800 ;
        RECT 84.600 95.200 84.900 108.800 ;
        RECT 85.400 103.100 85.800 108.900 ;
        RECT 87.000 108.800 87.400 109.200 ;
        RECT 89.400 108.800 89.800 109.200 ;
        RECT 89.400 106.300 89.700 108.800 ;
        RECT 89.400 105.800 89.800 106.300 ;
        RECT 90.200 103.100 90.600 108.900 ;
        RECT 91.000 107.200 91.300 112.800 ;
        RECT 91.800 111.800 92.200 112.200 ;
        RECT 95.000 111.800 95.400 112.200 ;
        RECT 97.400 112.100 97.800 117.900 ;
        RECT 98.200 113.800 98.600 114.200 ;
        RECT 98.200 113.200 98.500 113.800 ;
        RECT 98.200 112.800 98.600 113.200 ;
        RECT 91.800 109.200 92.100 111.800 ;
        RECT 95.000 111.200 95.300 111.800 ;
        RECT 95.000 110.800 95.400 111.200 ;
        RECT 94.200 109.800 94.600 110.200 ;
        RECT 94.200 109.200 94.500 109.800 ;
        RECT 95.000 109.200 95.300 110.800 ;
        RECT 91.800 108.800 92.200 109.200 ;
        RECT 94.200 108.800 94.600 109.200 ;
        RECT 95.000 108.800 95.400 109.200 ;
        RECT 91.000 106.800 91.400 107.200 ;
        RECT 87.000 98.100 87.400 98.200 ;
        RECT 87.800 98.100 88.200 98.200 ;
        RECT 87.000 97.800 88.200 98.100 ;
        RECT 73.400 94.800 73.800 95.200 ;
        RECT 74.200 94.800 74.600 95.200 ;
        RECT 77.400 94.800 77.800 95.200 ;
        RECT 80.600 94.800 81.000 95.200 ;
        RECT 81.400 94.800 81.800 95.200 ;
        RECT 83.800 94.800 84.200 95.200 ;
        RECT 84.600 94.800 85.000 95.200 ;
        RECT 87.000 94.800 87.400 95.200 ;
        RECT 72.600 88.800 73.000 89.200 ;
        RECT 71.800 84.800 72.200 85.200 ;
        RECT 71.800 82.200 72.100 84.800 ;
        RECT 71.800 81.800 72.200 82.200 ;
        RECT 73.400 76.100 73.700 94.800 ;
        RECT 74.200 89.200 74.500 94.800 ;
        RECT 74.200 88.800 74.600 89.200 ;
        RECT 76.600 83.100 77.000 88.900 ;
        RECT 72.600 75.800 73.700 76.100 ;
        RECT 70.200 74.800 70.600 75.200 ;
        RECT 70.200 72.200 70.500 74.800 ;
        RECT 70.200 71.800 70.600 72.200 ;
        RECT 62.200 67.800 62.600 68.200 ;
        RECT 63.800 67.800 64.200 68.200 ;
        RECT 59.800 66.800 60.200 67.200 ;
        RECT 59.000 65.800 59.400 66.200 ;
        RECT 59.800 66.100 60.200 66.200 ;
        RECT 60.600 66.100 61.000 66.200 ;
        RECT 59.800 65.800 61.000 66.100 ;
        RECT 59.000 65.200 59.300 65.800 ;
        RECT 53.400 64.800 53.800 65.200 ;
        RECT 57.400 64.800 57.800 65.200 ;
        RECT 59.000 64.800 59.400 65.200 ;
        RECT 48.600 61.800 49.000 62.200 ;
        RECT 60.600 61.800 61.000 62.200 ;
        RECT 44.600 55.800 45.000 56.200 ;
        RECT 45.400 55.800 45.800 56.200 ;
        RECT 44.600 55.200 44.900 55.800 ;
        RECT 44.600 54.800 45.000 55.200 ;
        RECT 35.800 52.800 36.200 53.200 ;
        RECT 42.200 52.800 42.600 53.200 ;
        RECT 43.000 52.800 43.400 53.200 ;
        RECT 27.800 49.800 28.200 50.200 ;
        RECT 27.000 47.800 27.400 48.200 ;
        RECT 27.800 46.200 28.100 49.800 ;
        RECT 30.200 49.200 30.500 52.800 ;
        RECT 32.600 51.800 33.000 52.200 ;
        RECT 28.600 48.800 29.000 49.200 ;
        RECT 30.200 48.800 30.600 49.200 ;
        RECT 27.800 45.800 28.200 46.200 ;
        RECT 22.200 39.800 22.600 40.200 ;
        RECT 14.200 34.800 14.600 35.200 ;
        RECT 17.400 32.100 17.800 37.900 ;
        RECT 19.000 33.100 19.400 35.900 ;
        RECT 19.800 33.100 20.200 35.900 ;
        RECT 21.400 32.100 21.800 37.900 ;
        RECT 22.200 35.100 22.500 39.800 ;
        RECT 28.600 39.200 28.900 48.800 ;
        RECT 30.200 47.800 30.600 48.200 ;
        RECT 30.200 46.200 30.500 47.800 ;
        RECT 30.200 45.800 30.600 46.200 ;
        RECT 31.000 43.100 31.400 48.900 ;
        RECT 32.600 47.200 32.900 51.800 ;
        RECT 43.000 50.200 43.300 52.800 ;
        RECT 33.400 49.800 33.800 50.200 ;
        RECT 38.200 49.800 38.600 50.200 ;
        RECT 40.600 49.800 41.000 50.200 ;
        RECT 43.000 49.800 43.400 50.200 ;
        RECT 33.400 49.200 33.700 49.800 ;
        RECT 38.200 49.200 38.500 49.800 ;
        RECT 33.400 48.800 33.800 49.200 ;
        RECT 38.200 48.800 38.600 49.200 ;
        RECT 39.000 48.800 39.400 49.200 ;
        RECT 39.000 48.200 39.300 48.800 ;
        RECT 39.000 47.800 39.400 48.200 ;
        RECT 40.600 47.200 40.900 49.800 ;
        RECT 42.200 49.100 42.600 49.200 ;
        RECT 43.000 49.100 43.400 49.200 ;
        RECT 42.200 48.800 43.400 49.100 ;
        RECT 41.400 47.500 41.800 47.900 ;
        RECT 44.500 47.800 44.900 47.900 ;
        RECT 42.100 47.500 44.900 47.800 ;
        RECT 32.600 46.800 33.000 47.200 ;
        RECT 37.400 47.100 37.800 47.200 ;
        RECT 38.200 47.100 38.600 47.200 ;
        RECT 37.400 46.800 38.600 47.100 ;
        RECT 40.600 46.800 41.000 47.200 ;
        RECT 41.400 47.100 41.700 47.500 ;
        RECT 42.100 47.400 42.500 47.500 ;
        RECT 43.800 47.400 44.200 47.500 ;
        RECT 41.400 46.800 44.200 47.100 ;
        RECT 35.800 42.800 36.200 43.200 ;
        RECT 28.600 38.800 29.000 39.200 ;
        RECT 22.200 34.700 22.600 35.100 ;
        RECT 23.800 34.100 24.200 34.200 ;
        RECT 24.600 34.100 25.000 34.200 ;
        RECT 23.800 33.800 25.000 34.100 ;
        RECT 11.000 29.800 11.400 30.200 ;
        RECT 8.600 28.800 9.700 29.100 ;
        RECT 8.600 25.100 9.000 27.900 ;
        RECT 9.400 27.200 9.700 28.800 ;
        RECT 9.400 26.800 9.800 27.200 ;
        RECT 7.000 24.100 7.400 24.200 ;
        RECT 7.800 24.100 8.200 24.200 ;
        RECT 7.000 23.800 8.200 24.100 ;
        RECT 10.200 23.100 10.600 28.900 ;
        RECT 0.600 11.800 1.000 12.200 ;
        RECT 3.000 12.100 3.400 12.200 ;
        RECT 3.800 12.100 4.200 12.200 ;
        RECT 5.400 12.100 5.800 17.900 ;
        RECT 8.600 14.800 9.000 15.200 ;
        RECT 3.000 11.800 4.200 12.100 ;
        RECT 0.600 8.200 0.900 11.800 ;
        RECT 7.000 10.800 7.400 11.200 ;
        RECT 7.000 8.200 7.300 10.800 ;
        RECT 0.600 7.800 1.000 8.200 ;
        RECT 7.000 7.800 7.400 8.200 ;
        RECT 8.600 7.200 8.900 14.800 ;
        RECT 10.200 12.100 10.600 17.900 ;
        RECT 11.000 16.200 11.300 29.800 ;
        RECT 14.200 27.800 14.600 28.200 ;
        RECT 14.200 27.200 14.500 27.800 ;
        RECT 14.200 26.800 14.600 27.200 ;
        RECT 11.800 26.100 12.200 26.200 ;
        RECT 12.600 26.100 13.000 26.200 ;
        RECT 11.800 25.800 13.000 26.100 ;
        RECT 15.000 23.100 15.400 28.900 ;
        RECT 18.200 25.100 18.600 27.900 ;
        RECT 19.800 23.100 20.200 28.900 ;
        RECT 20.600 25.900 21.000 26.300 ;
        RECT 23.800 26.200 24.100 33.800 ;
        RECT 26.200 32.100 26.600 37.900 ;
        RECT 28.600 36.200 28.900 38.800 ;
        RECT 28.600 35.800 29.000 36.200 ;
        RECT 29.400 32.100 29.800 32.200 ;
        RECT 30.200 32.100 30.600 32.200 ;
        RECT 31.800 32.100 32.200 37.900 ;
        RECT 35.800 35.100 36.100 42.800 ;
        RECT 40.600 39.200 40.900 46.800 ;
        RECT 41.400 45.100 41.700 46.800 ;
        RECT 42.200 46.100 42.600 46.200 ;
        RECT 43.900 46.100 44.200 46.800 ;
        RECT 42.200 45.800 43.300 46.100 ;
        RECT 41.400 44.700 41.800 45.100 ;
        RECT 43.000 39.200 43.300 45.800 ;
        RECT 43.900 45.700 44.300 46.100 ;
        RECT 44.600 45.100 44.900 47.500 ;
        RECT 45.400 47.200 45.700 55.800 ;
        RECT 48.600 55.200 48.900 61.800 ;
        RECT 51.000 57.800 51.400 58.200 ;
        RECT 51.000 56.200 51.300 57.800 ;
        RECT 51.800 56.800 52.200 57.200 ;
        RECT 51.800 56.200 52.100 56.800 ;
        RECT 49.400 55.800 49.800 56.200 ;
        RECT 51.000 55.800 51.400 56.200 ;
        RECT 51.800 55.800 52.200 56.200 ;
        RECT 48.600 54.800 49.000 55.200 ;
        RECT 49.400 54.200 49.700 55.800 ;
        RECT 51.000 54.800 51.400 55.200 ;
        RECT 49.400 53.800 49.800 54.200 ;
        RECT 47.800 52.800 48.200 53.200 ;
        RECT 47.800 49.200 48.100 52.800 ;
        RECT 47.800 49.100 48.200 49.200 ;
        RECT 48.600 49.100 49.000 49.200 ;
        RECT 47.800 48.800 49.000 49.100 ;
        RECT 45.400 46.800 45.800 47.200 ;
        RECT 44.500 44.700 44.900 45.100 ;
        RECT 50.200 43.100 50.600 48.900 ;
        RECT 47.800 41.800 48.200 42.200 ;
        RECT 40.600 38.800 41.000 39.200 ;
        RECT 43.000 38.800 43.400 39.200 ;
        RECT 35.800 34.700 36.200 35.100 ;
        RECT 35.800 34.200 36.100 34.700 ;
        RECT 32.600 33.800 33.000 34.200 ;
        RECT 35.800 33.800 36.200 34.200 ;
        RECT 32.600 33.200 32.900 33.800 ;
        RECT 32.600 32.800 33.000 33.200 ;
        RECT 35.800 32.800 36.200 33.200 ;
        RECT 29.400 31.800 30.600 32.100 ;
        RECT 20.600 25.200 20.900 25.900 ;
        RECT 23.800 25.800 24.200 26.200 ;
        RECT 20.600 24.800 21.000 25.200 ;
        RECT 17.400 22.100 17.800 22.200 ;
        RECT 18.200 22.100 18.600 22.200 ;
        RECT 17.400 21.800 18.600 22.100 ;
        RECT 11.000 15.800 11.400 16.200 ;
        RECT 11.000 14.200 11.300 15.800 ;
        RECT 11.000 13.800 11.400 14.200 ;
        RECT 11.800 13.100 12.200 15.900 ;
        RECT 12.600 14.800 13.000 15.200 ;
        RECT 12.600 10.200 12.900 14.800 ;
        RECT 14.200 12.800 14.600 13.200 ;
        RECT 15.000 13.100 15.400 15.900 ;
        RECT 14.200 12.200 14.500 12.800 ;
        RECT 13.400 11.800 13.800 12.200 ;
        RECT 14.200 11.800 14.600 12.200 ;
        RECT 16.600 12.100 17.000 17.900 ;
        RECT 17.400 14.700 17.800 15.100 ;
        RECT 17.400 14.200 17.700 14.700 ;
        RECT 17.400 13.800 17.800 14.200 ;
        RECT 13.400 11.200 13.700 11.800 ;
        RECT 13.400 10.800 13.800 11.200 ;
        RECT 12.600 9.800 13.000 10.200 ;
        RECT 11.800 9.100 12.200 9.200 ;
        RECT 12.600 9.100 13.000 9.200 ;
        RECT 11.800 8.800 13.000 9.100 ;
        RECT 12.600 8.100 13.000 8.200 ;
        RECT 13.400 8.100 13.800 8.200 ;
        RECT 12.600 7.800 13.800 8.100 ;
        RECT 15.800 7.800 16.200 8.200 ;
        RECT 16.600 8.100 17.000 8.200 ;
        RECT 17.400 8.100 17.800 8.200 ;
        RECT 16.600 7.800 17.800 8.100 ;
        RECT 15.800 7.200 16.100 7.800 ;
        RECT 18.200 7.200 18.500 21.800 ;
        RECT 20.600 16.800 21.000 17.200 ;
        RECT 20.600 15.200 20.900 16.800 ;
        RECT 19.000 14.800 19.400 15.200 ;
        RECT 20.600 14.800 21.000 15.200 ;
        RECT 19.000 9.200 19.300 14.800 ;
        RECT 21.400 12.100 21.800 17.900 ;
        RECT 23.800 17.200 24.100 25.800 ;
        RECT 24.600 23.100 25.000 28.900 ;
        RECT 27.800 25.100 28.200 27.900 ;
        RECT 28.600 27.800 29.000 28.200 ;
        RECT 28.600 27.200 28.900 27.800 ;
        RECT 28.600 26.800 29.000 27.200 ;
        RECT 25.400 22.800 25.800 23.200 ;
        RECT 29.400 23.100 29.800 28.900 ;
        RECT 30.200 25.900 30.600 26.300 ;
        RECT 30.200 23.200 30.500 25.900 ;
        RECT 30.200 22.800 30.600 23.200 ;
        RECT 34.200 23.100 34.600 28.900 ;
        RECT 35.000 28.800 35.400 29.200 ;
        RECT 25.400 19.200 25.700 22.800 ;
        RECT 26.200 22.100 26.600 22.200 ;
        RECT 27.000 22.100 27.400 22.200 ;
        RECT 26.200 21.800 27.400 22.100 ;
        RECT 25.400 18.800 25.800 19.200 ;
        RECT 35.000 17.200 35.300 28.800 ;
        RECT 35.800 27.100 36.100 32.800 ;
        RECT 36.600 32.100 37.000 37.900 ;
        RECT 47.800 36.200 48.100 41.800 ;
        RECT 38.200 33.100 38.600 35.900 ;
        RECT 39.000 35.800 39.400 36.200 ;
        RECT 47.800 35.800 48.200 36.200 ;
        RECT 50.200 35.800 50.600 36.200 ;
        RECT 39.000 34.200 39.300 35.800 ;
        RECT 39.800 35.100 40.200 35.200 ;
        RECT 40.600 35.100 41.000 35.200 ;
        RECT 39.800 34.800 41.000 35.100 ;
        RECT 43.000 34.800 43.400 35.200 ;
        RECT 44.600 35.100 45.000 35.200 ;
        RECT 45.400 35.100 45.800 35.200 ;
        RECT 44.600 34.800 45.800 35.100 ;
        RECT 49.400 34.800 49.800 35.200 ;
        RECT 39.000 33.800 39.400 34.200 ;
        RECT 42.200 33.800 42.600 34.200 ;
        RECT 38.200 30.800 38.600 31.200 ;
        RECT 38.200 29.200 38.500 30.800 ;
        RECT 36.600 28.800 37.000 29.200 ;
        RECT 38.200 28.800 38.600 29.200 ;
        RECT 36.600 28.200 36.900 28.800 ;
        RECT 39.000 28.200 39.300 33.800 ;
        RECT 36.600 27.800 37.000 28.200 ;
        RECT 39.000 27.800 39.400 28.200 ;
        RECT 35.800 26.800 36.900 27.100 ;
        RECT 36.600 17.200 36.900 26.800 ;
        RECT 37.400 26.100 37.800 26.200 ;
        RECT 38.200 26.100 38.600 26.200 ;
        RECT 37.400 25.800 38.600 26.100 ;
        RECT 39.800 25.100 40.200 27.900 ;
        RECT 40.600 27.800 41.000 28.200 ;
        RECT 40.600 27.200 40.900 27.800 ;
        RECT 40.600 26.800 41.000 27.200 ;
        RECT 40.600 22.800 41.000 23.200 ;
        RECT 41.400 23.100 41.800 28.900 ;
        RECT 42.200 26.300 42.500 33.800 ;
        RECT 43.000 31.200 43.300 34.800 ;
        RECT 49.400 34.200 49.700 34.800 ;
        RECT 50.200 34.200 50.500 35.800 ;
        RECT 51.000 35.200 51.300 54.800 ;
        RECT 54.200 52.100 54.600 57.900 ;
        RECT 57.400 55.000 57.800 55.100 ;
        RECT 58.200 55.000 58.600 55.100 ;
        RECT 57.400 54.700 58.600 55.000 ;
        RECT 57.400 53.800 57.800 54.200 ;
        RECT 58.200 53.800 58.600 54.200 ;
        RECT 57.400 53.200 57.700 53.800 ;
        RECT 57.400 52.800 57.800 53.200 ;
        RECT 53.400 46.200 53.800 46.300 ;
        RECT 54.200 46.200 54.600 46.300 ;
        RECT 53.400 45.900 54.600 46.200 ;
        RECT 55.000 43.100 55.400 48.900 ;
        RECT 55.800 47.800 56.200 48.200 ;
        RECT 55.800 47.200 56.100 47.800 ;
        RECT 55.800 46.800 56.200 47.200 ;
        RECT 56.600 45.100 57.000 47.900 ;
        RECT 52.600 39.100 53.000 39.200 ;
        RECT 53.400 39.100 53.800 39.200 ;
        RECT 52.600 38.800 53.800 39.100 ;
        RECT 51.000 34.800 51.400 35.200 ;
        RECT 51.800 35.100 52.200 35.200 ;
        RECT 52.600 35.100 53.000 35.200 ;
        RECT 51.800 34.800 53.000 35.100 ;
        RECT 51.000 34.200 51.300 34.800 ;
        RECT 49.400 33.800 49.800 34.200 ;
        RECT 50.200 33.800 50.600 34.200 ;
        RECT 51.000 33.800 51.400 34.200 ;
        RECT 54.200 33.800 54.600 34.200 ;
        RECT 50.200 33.200 50.500 33.800 ;
        RECT 50.200 32.800 50.600 33.200 ;
        RECT 52.600 33.100 53.000 33.200 ;
        RECT 53.400 33.100 53.800 33.200 ;
        RECT 52.600 32.800 53.800 33.100 ;
        RECT 43.000 30.800 43.400 31.200 ;
        RECT 54.200 29.200 54.500 33.800 ;
        RECT 55.800 32.100 56.200 37.900 ;
        RECT 57.400 35.200 57.700 52.800 ;
        RECT 58.200 48.200 58.500 53.800 ;
        RECT 59.000 52.100 59.400 57.900 ;
        RECT 60.600 57.100 60.900 61.800 ;
        RECT 59.800 56.800 60.900 57.100 ;
        RECT 61.400 56.800 61.800 57.200 ;
        RECT 58.200 47.800 58.600 48.200 ;
        RECT 58.200 47.200 58.500 47.800 ;
        RECT 58.200 46.800 58.600 47.200 ;
        RECT 57.400 34.800 57.800 35.200 ;
        RECT 59.800 35.100 60.100 56.800 ;
        RECT 61.400 56.200 61.700 56.800 ;
        RECT 60.600 53.100 61.000 55.900 ;
        RECT 61.400 55.800 61.800 56.200 ;
        RECT 63.800 52.100 64.200 57.900 ;
        RECT 64.600 55.200 64.900 71.800 ;
        RECT 67.000 70.200 67.300 71.800 ;
        RECT 67.000 69.800 67.400 70.200 ;
        RECT 65.400 63.100 65.800 68.900 ;
        RECT 69.400 66.800 69.800 67.200 ;
        RECT 69.400 66.300 69.700 66.800 ;
        RECT 69.400 65.900 69.800 66.300 ;
        RECT 70.200 63.100 70.600 68.900 ;
        RECT 71.000 67.800 71.400 68.200 ;
        RECT 71.000 67.200 71.300 67.800 ;
        RECT 71.000 66.800 71.400 67.200 ;
        RECT 71.800 65.100 72.200 67.900 ;
        RECT 72.600 66.200 72.900 75.800 ;
        RECT 73.400 74.700 73.800 75.100 ;
        RECT 73.400 73.200 73.700 74.700 ;
        RECT 73.400 72.800 73.800 73.200 ;
        RECT 73.400 67.200 73.700 72.800 ;
        RECT 74.200 72.100 74.600 77.900 ;
        RECT 77.400 76.200 77.700 94.800 ;
        RECT 79.800 93.100 80.200 93.200 ;
        RECT 80.600 93.100 81.000 93.200 ;
        RECT 79.800 92.800 81.000 93.100 ;
        RECT 81.400 92.200 81.700 94.800 ;
        RECT 79.000 91.800 79.400 92.200 ;
        RECT 81.400 91.800 81.800 92.200 ;
        RECT 79.000 86.200 79.300 91.800 ;
        RECT 84.600 89.200 84.900 94.800 ;
        RECT 87.000 94.200 87.300 94.800 ;
        RECT 87.000 93.800 87.400 94.200 ;
        RECT 87.000 93.100 87.400 93.200 ;
        RECT 87.800 93.100 88.200 93.200 ;
        RECT 87.000 92.800 88.200 93.100 ;
        RECT 87.800 91.800 88.200 92.200 ;
        RECT 90.200 92.100 90.600 97.900 ;
        RECT 91.000 95.200 91.300 106.800 ;
        RECT 91.800 105.100 92.200 107.900 ;
        RECT 96.600 103.100 97.000 108.900 ;
        RECT 99.000 107.200 99.300 126.800 ;
        RECT 99.800 125.100 100.200 127.900 ;
        RECT 100.600 125.200 100.900 134.800 ;
        RECT 103.000 129.200 103.300 147.800 ;
        RECT 103.800 139.200 104.100 147.800 ;
        RECT 106.200 143.100 106.600 148.900 ;
        RECT 107.000 145.800 107.400 146.200 ;
        RECT 107.000 145.200 107.300 145.800 ;
        RECT 107.000 144.800 107.400 145.200 ;
        RECT 108.600 139.200 108.900 152.800 ;
        RECT 110.200 151.200 110.500 154.800 ;
        RECT 110.200 150.800 110.600 151.200 ;
        RECT 113.400 149.200 113.700 154.800 ;
        RECT 110.200 146.800 110.600 147.200 ;
        RECT 110.200 146.300 110.500 146.800 ;
        RECT 110.200 145.900 110.600 146.300 ;
        RECT 111.000 143.100 111.400 148.900 ;
        RECT 113.400 148.800 113.800 149.200 ;
        RECT 112.600 145.100 113.000 147.900 ;
        RECT 113.400 141.800 113.800 142.200 ;
        RECT 103.800 138.800 104.200 139.200 ;
        RECT 108.600 138.800 109.000 139.200 ;
        RECT 113.400 136.200 113.700 141.800 ;
        RECT 115.000 139.200 115.300 154.800 ;
        RECT 121.400 154.100 121.800 154.200 ;
        RECT 122.200 154.100 122.600 154.200 ;
        RECT 121.400 153.800 122.600 154.100 ;
        RECT 125.400 153.800 125.800 154.200 ;
        RECT 117.400 152.800 117.800 153.200 ;
        RECT 119.000 153.100 119.400 153.200 ;
        RECT 119.800 153.100 120.200 153.200 ;
        RECT 119.000 152.800 120.200 153.100 ;
        RECT 115.800 143.100 116.200 148.900 ;
        RECT 117.400 148.200 117.700 152.800 ;
        RECT 119.800 152.200 120.100 152.800 ;
        RECT 125.400 152.200 125.700 153.800 ;
        RECT 127.800 153.200 128.100 154.800 ;
        RECT 130.200 154.200 130.500 154.800 ;
        RECT 130.200 153.800 130.600 154.200 ;
        RECT 127.800 152.800 128.200 153.200 ;
        RECT 129.400 152.800 129.800 153.200 ;
        RECT 119.800 151.800 120.200 152.200 ;
        RECT 125.400 151.800 125.800 152.200 ;
        RECT 127.000 150.800 127.400 151.200 ;
        RECT 117.400 147.800 117.800 148.200 ;
        RECT 119.000 146.200 119.400 146.300 ;
        RECT 119.800 146.200 120.200 146.300 ;
        RECT 119.000 145.900 120.200 146.200 ;
        RECT 119.800 142.800 120.200 143.200 ;
        RECT 120.600 143.100 121.000 148.900 ;
        RECT 121.400 147.800 121.800 148.200 ;
        RECT 123.000 148.100 123.400 148.200 ;
        RECT 123.800 148.100 124.200 148.200 ;
        RECT 121.400 147.200 121.700 147.800 ;
        RECT 121.400 146.800 121.800 147.200 ;
        RECT 122.200 145.100 122.600 147.900 ;
        RECT 123.000 147.800 124.200 148.100 ;
        RECT 124.600 148.100 125.000 148.200 ;
        RECT 124.600 147.800 125.700 148.100 ;
        RECT 124.600 147.200 124.900 147.800 ;
        RECT 125.400 147.200 125.700 147.800 ;
        RECT 126.200 147.800 126.600 148.200 ;
        RECT 124.600 146.800 125.000 147.200 ;
        RECT 125.400 146.800 125.800 147.200 ;
        RECT 123.000 146.100 123.400 146.200 ;
        RECT 123.000 145.800 124.100 146.100 ;
        RECT 119.800 139.200 120.100 142.800 ;
        RECT 123.800 139.200 124.100 145.800 ;
        RECT 115.000 138.800 115.400 139.200 ;
        RECT 119.800 138.800 120.200 139.200 ;
        RECT 123.800 138.800 124.200 139.200 ;
        RECT 113.400 135.800 113.800 136.200 ;
        RECT 125.400 135.800 125.800 136.200 ;
        RECT 125.400 135.200 125.700 135.800 ;
        RECT 126.200 135.200 126.500 147.800 ;
        RECT 127.000 135.200 127.300 150.800 ;
        RECT 127.800 143.200 128.100 152.800 ;
        RECT 127.800 142.800 128.200 143.200 ;
        RECT 127.800 141.800 128.200 142.200 ;
        RECT 127.800 135.200 128.100 141.800 ;
        RECT 129.400 139.200 129.700 152.800 ;
        RECT 129.400 138.800 129.800 139.200 ;
        RECT 131.000 138.200 131.300 157.800 ;
        RECT 132.600 154.800 133.000 155.200 ;
        RECT 134.200 154.800 134.600 155.200 ;
        RECT 132.600 153.200 132.900 154.800 ;
        RECT 134.200 154.200 134.500 154.800 ;
        RECT 134.200 153.800 134.600 154.200 ;
        RECT 132.600 152.800 133.000 153.200 ;
        RECT 134.200 152.800 134.600 153.200 ;
        RECT 132.600 151.800 133.000 152.200 ;
        RECT 132.600 149.200 132.900 151.800 ;
        RECT 132.600 148.800 133.000 149.200 ;
        RECT 134.200 147.200 134.500 152.800 ;
        RECT 135.000 151.800 135.400 152.200 ;
        RECT 137.400 152.100 137.800 157.900 ;
        RECT 138.200 155.200 138.500 166.800 ;
        RECT 139.000 166.200 139.300 166.800 ;
        RECT 139.000 165.800 139.400 166.200 ;
        RECT 142.200 163.100 142.600 168.900 ;
        RECT 144.600 168.100 145.000 168.200 ;
        RECT 145.400 168.100 145.800 168.200 ;
        RECT 144.600 167.800 145.800 168.100 ;
        RECT 151.000 167.800 151.400 168.200 ;
        RECT 151.000 167.200 151.300 167.800 ;
        RECT 145.400 166.800 145.800 167.200 ;
        RECT 147.000 166.800 147.400 167.200 ;
        RECT 151.000 166.800 151.400 167.200 ;
        RECT 145.400 166.200 145.700 166.800 ;
        RECT 147.000 166.200 147.300 166.800 ;
        RECT 144.600 165.800 145.000 166.200 ;
        RECT 145.400 165.800 145.800 166.200 ;
        RECT 147.000 165.800 147.400 166.200 ;
        RECT 149.400 165.800 149.800 166.200 ;
        RECT 150.200 166.100 150.600 166.200 ;
        RECT 151.000 166.100 151.400 166.200 ;
        RECT 150.200 165.800 151.400 166.100 ;
        RECT 144.600 162.200 144.900 165.800 ;
        RECT 149.400 165.100 149.700 165.800 ;
        RECT 149.400 164.800 150.500 165.100 ;
        RECT 144.600 161.800 145.000 162.200 ;
        RECT 144.600 158.200 144.900 161.800 ;
        RECT 147.800 158.800 148.200 159.200 ;
        RECT 138.200 154.800 138.600 155.200 ;
        RECT 139.000 154.800 139.400 155.200 ;
        RECT 139.800 155.100 140.200 155.200 ;
        RECT 140.600 155.100 141.000 155.200 ;
        RECT 139.800 154.800 141.000 155.100 ;
        RECT 138.200 153.200 138.500 154.800 ;
        RECT 138.200 152.800 138.600 153.200 ;
        RECT 135.000 151.200 135.300 151.800 ;
        RECT 135.000 150.800 135.400 151.200 ;
        RECT 134.200 146.800 134.600 147.200 ;
        RECT 135.000 143.100 135.400 148.900 ;
        RECT 139.000 146.300 139.300 154.800 ;
        RECT 142.200 152.100 142.600 157.900 ;
        RECT 144.600 157.800 145.000 158.200 ;
        RECT 143.800 153.100 144.200 155.900 ;
        RECT 146.200 155.800 146.600 156.200 ;
        RECT 146.200 155.200 146.500 155.800 ;
        RECT 147.800 155.200 148.100 158.800 ;
        RECT 150.200 155.200 150.500 164.800 ;
        RECT 156.600 163.100 157.000 168.900 ;
        RECT 159.800 166.800 160.200 167.200 ;
        RECT 160.600 166.800 161.000 167.200 ;
        RECT 159.800 166.200 160.100 166.800 ;
        RECT 159.800 165.800 160.200 166.200 ;
        RECT 154.200 162.100 154.600 162.200 ;
        RECT 155.000 162.100 155.400 162.200 ;
        RECT 154.200 161.800 155.400 162.100 ;
        RECT 151.000 155.800 151.400 156.200 ;
        RECT 151.000 155.200 151.300 155.800 ;
        RECT 144.600 154.800 145.000 155.200 ;
        RECT 145.400 154.800 145.800 155.200 ;
        RECT 146.200 154.800 146.600 155.200 ;
        RECT 147.800 154.800 148.200 155.200 ;
        RECT 148.600 154.800 149.000 155.200 ;
        RECT 150.200 154.800 150.600 155.200 ;
        RECT 151.000 154.800 151.400 155.200 ;
        RECT 144.600 154.200 144.900 154.800 ;
        RECT 144.600 153.800 145.000 154.200 ;
        RECT 145.400 149.200 145.700 154.800 ;
        RECT 135.800 145.800 136.200 146.200 ;
        RECT 139.000 145.900 139.400 146.300 ;
        RECT 135.800 145.200 136.100 145.800 ;
        RECT 135.800 144.800 136.200 145.200 ;
        RECT 139.800 143.100 140.200 148.900 ;
        RECT 145.400 148.800 145.800 149.200 ;
        RECT 147.000 149.100 147.400 149.200 ;
        RECT 147.800 149.100 148.200 149.200 ;
        RECT 147.000 148.800 148.200 149.100 ;
        RECT 148.600 148.200 148.900 154.800 ;
        RECT 152.600 153.800 153.000 154.200 ;
        RECT 152.600 153.200 152.900 153.800 ;
        RECT 151.000 153.100 151.400 153.200 ;
        RECT 151.800 153.100 152.200 153.200 ;
        RECT 151.000 152.800 152.200 153.100 ;
        RECT 152.600 152.800 153.000 153.200 ;
        RECT 153.400 153.100 153.800 155.900 ;
        RECT 154.200 154.800 154.600 155.200 ;
        RECT 154.200 154.200 154.500 154.800 ;
        RECT 154.200 153.800 154.600 154.200 ;
        RECT 154.200 152.800 154.600 153.200 ;
        RECT 141.400 145.100 141.800 147.900 ;
        RECT 148.600 147.800 149.000 148.200 ;
        RECT 148.600 146.200 148.900 147.800 ;
        RECT 148.600 145.800 149.000 146.200 ;
        RECT 151.000 145.100 151.400 147.900 ;
        RECT 151.800 146.800 152.200 147.200 ;
        RECT 151.800 145.200 152.100 146.800 ;
        RECT 151.800 144.800 152.200 145.200 ;
        RECT 152.600 143.100 153.000 148.900 ;
        RECT 154.200 146.200 154.500 152.800 ;
        RECT 155.000 152.100 155.400 157.900 ;
        RECT 156.600 154.800 157.000 155.200 ;
        RECT 156.600 153.200 156.900 154.800 ;
        RECT 156.600 152.800 157.000 153.200 ;
        RECT 159.800 152.100 160.200 157.900 ;
        RECT 160.600 157.200 160.900 166.800 ;
        RECT 161.400 163.100 161.800 168.900 ;
        RECT 163.000 165.100 163.400 167.900 ;
        RECT 163.800 165.100 164.200 167.900 ;
        RECT 163.000 163.800 163.400 164.200 ;
        RECT 161.400 159.100 161.800 159.200 ;
        RECT 162.200 159.100 162.600 159.200 ;
        RECT 161.400 158.800 162.600 159.100 ;
        RECT 163.000 158.100 163.300 163.800 ;
        RECT 165.400 163.100 165.800 168.900 ;
        RECT 167.000 165.800 167.400 166.200 ;
        RECT 169.400 165.800 169.800 166.200 ;
        RECT 167.000 159.200 167.300 165.800 ;
        RECT 169.400 165.200 169.700 165.800 ;
        RECT 169.400 164.800 169.800 165.200 ;
        RECT 170.200 163.100 170.600 168.900 ;
        RECT 178.200 163.100 178.600 168.900 ;
        RECT 179.000 166.100 179.400 166.200 ;
        RECT 179.800 166.100 180.200 166.200 ;
        RECT 179.000 165.800 180.200 166.100 ;
        RECT 181.400 165.800 181.800 166.200 ;
        RECT 172.600 161.800 173.000 162.200 ;
        RECT 175.800 161.800 176.200 162.200 ;
        RECT 167.000 158.800 167.400 159.200 ;
        RECT 162.200 157.800 163.300 158.100 ;
        RECT 160.600 156.800 161.000 157.200 ;
        RECT 160.600 152.800 161.000 153.200 ;
        RECT 159.800 149.100 160.200 149.200 ;
        RECT 160.600 149.100 160.900 152.800 ;
        RECT 154.200 145.800 154.600 146.200 ;
        RECT 157.400 143.100 157.800 148.900 ;
        RECT 159.800 148.800 160.900 149.100 ;
        RECT 162.200 149.200 162.500 157.800 ;
        RECT 171.800 154.800 172.200 155.200 ;
        RECT 166.200 153.800 166.600 154.200 ;
        RECT 166.200 153.200 166.500 153.800 ;
        RECT 171.800 153.200 172.100 154.800 ;
        RECT 166.200 152.800 166.600 153.200 ;
        RECT 171.800 153.100 172.200 153.200 ;
        RECT 172.600 153.100 172.900 161.800 ;
        RECT 175.800 158.200 176.100 161.800 ;
        RECT 181.400 159.200 181.700 165.800 ;
        RECT 183.000 163.100 183.400 168.900 ;
        RECT 183.800 166.800 184.200 167.200 ;
        RECT 181.400 158.800 181.800 159.200 ;
        RECT 175.800 157.800 176.200 158.200 ;
        RECT 175.800 155.200 176.100 157.800 ;
        RECT 181.400 155.200 181.700 158.800 ;
        RECT 171.800 152.800 172.900 153.100 ;
        RECT 173.400 154.800 173.800 155.200 ;
        RECT 174.200 154.800 174.600 155.200 ;
        RECT 175.800 154.800 176.200 155.200 ;
        RECT 177.400 154.800 177.800 155.200 ;
        RECT 180.600 154.800 181.000 155.200 ;
        RECT 181.400 154.800 181.800 155.200 ;
        RECT 163.000 151.800 163.400 152.200 ;
        RECT 162.200 148.800 162.600 149.200 ;
        RECT 163.000 148.200 163.300 151.800 ;
        RECT 171.800 148.800 172.200 149.200 ;
        RECT 171.800 148.200 172.100 148.800 ;
        RECT 163.000 147.800 163.400 148.200 ;
        RECT 167.000 147.800 167.400 148.200 ;
        RECT 171.800 147.800 172.200 148.200 ;
        RECT 167.000 147.200 167.300 147.800 ;
        RECT 160.600 147.100 161.000 147.200 ;
        RECT 161.400 147.100 161.800 147.200 ;
        RECT 160.600 146.800 161.800 147.100 ;
        RECT 167.000 146.800 167.400 147.200 ;
        RECT 162.200 146.100 162.600 146.200 ;
        RECT 163.000 146.100 163.400 146.200 ;
        RECT 162.200 145.800 163.400 146.100 ;
        RECT 163.800 145.800 164.200 146.200 ;
        RECT 170.200 145.800 170.600 146.200 ;
        RECT 162.200 145.100 162.600 145.200 ;
        RECT 163.000 145.100 163.400 145.200 ;
        RECT 162.200 144.800 163.400 145.100 ;
        RECT 163.800 143.200 164.100 145.800 ;
        RECT 170.200 145.200 170.500 145.800 ;
        RECT 165.400 145.100 165.800 145.200 ;
        RECT 166.200 145.100 166.600 145.200 ;
        RECT 165.400 144.800 166.600 145.100 ;
        RECT 170.200 144.800 170.600 145.200 ;
        RECT 171.000 144.800 171.400 145.200 ;
        RECT 172.600 145.100 173.000 147.900 ;
        RECT 173.400 146.200 173.700 154.800 ;
        RECT 174.200 154.200 174.500 154.800 ;
        RECT 177.400 154.200 177.700 154.800 ;
        RECT 180.600 154.200 180.900 154.800 ;
        RECT 174.200 153.800 174.600 154.200 ;
        RECT 177.400 153.800 177.800 154.200 ;
        RECT 180.600 153.800 181.000 154.200 ;
        RECT 182.200 152.800 182.600 153.200 ;
        RECT 183.000 153.100 183.400 155.900 ;
        RECT 182.200 149.200 182.500 152.800 ;
        RECT 183.800 152.100 184.100 166.800 ;
        RECT 184.600 165.100 185.000 167.900 ;
        RECT 192.600 167.800 193.000 168.200 ;
        RECT 192.600 164.200 192.900 167.800 ;
        RECT 192.600 163.800 193.000 164.200 ;
        RECT 194.200 161.800 194.600 162.200 ;
        RECT 191.000 158.100 191.400 158.200 ;
        RECT 191.800 158.100 192.200 158.200 ;
        RECT 184.600 152.100 185.000 157.900 ;
        RECT 185.400 155.800 185.800 156.200 ;
        RECT 185.400 155.100 185.700 155.800 ;
        RECT 185.400 154.700 185.800 155.100 ;
        RECT 189.400 152.100 189.800 157.900 ;
        RECT 191.000 157.800 192.200 158.100 ;
        RECT 183.000 151.800 184.100 152.100 ;
        RECT 173.400 145.800 173.800 146.200 ;
        RECT 171.000 144.200 171.300 144.800 ;
        RECT 171.000 143.800 171.400 144.200 ;
        RECT 163.800 142.800 164.200 143.200 ;
        RECT 174.200 143.100 174.600 148.900 ;
        RECT 175.000 148.800 175.400 149.200 ;
        RECT 175.000 148.200 175.300 148.800 ;
        RECT 175.000 147.800 175.400 148.200 ;
        RECT 175.800 146.800 176.200 147.200 ;
        RECT 175.000 145.900 175.400 146.300 ;
        RECT 175.000 145.200 175.300 145.900 ;
        RECT 175.000 144.800 175.400 145.200 ;
        RECT 131.800 142.100 132.200 142.200 ;
        RECT 132.600 142.100 133.000 142.200 ;
        RECT 131.800 141.800 133.000 142.100 ;
        RECT 161.400 141.800 161.800 142.200 ;
        RECT 161.400 139.200 161.700 141.800 ;
        RECT 161.400 138.800 161.800 139.200 ;
        RECT 131.000 137.800 131.400 138.200 ;
        RECT 161.400 137.800 161.800 138.200 ;
        RECT 131.000 135.200 131.300 137.800 ;
        RECT 131.800 136.800 132.200 137.200 ;
        RECT 137.400 136.800 137.800 137.200 ;
        RECT 145.400 136.800 145.800 137.200 ;
        RECT 149.400 137.100 149.800 137.200 ;
        RECT 150.200 137.100 150.600 137.200 ;
        RECT 149.400 136.800 150.600 137.100 ;
        RECT 131.800 136.200 132.100 136.800 ;
        RECT 137.400 136.200 137.700 136.800 ;
        RECT 145.400 136.200 145.700 136.800 ;
        RECT 131.800 135.800 132.200 136.200 ;
        RECT 134.200 135.800 134.600 136.200 ;
        RECT 137.400 135.800 137.800 136.200 ;
        RECT 141.400 135.800 141.800 136.200 ;
        RECT 145.400 135.800 145.800 136.200 ;
        RECT 146.200 135.800 146.600 136.200 ;
        RECT 154.200 136.100 154.600 136.200 ;
        RECT 155.000 136.100 155.400 136.200 ;
        RECT 154.200 135.800 155.400 136.100 ;
        RECT 157.400 135.800 157.800 136.200 ;
        RECT 160.600 135.800 161.000 136.200 ;
        RECT 104.600 135.100 105.000 135.200 ;
        RECT 105.400 135.100 105.800 135.200 ;
        RECT 104.600 134.800 105.800 135.100 ;
        RECT 107.000 134.800 107.400 135.200 ;
        RECT 111.000 134.800 111.400 135.200 ;
        RECT 113.400 134.800 113.800 135.200 ;
        RECT 117.400 134.800 117.800 135.200 ;
        RECT 120.600 134.800 121.000 135.200 ;
        RECT 123.000 135.100 123.400 135.200 ;
        RECT 123.800 135.100 124.200 135.200 ;
        RECT 123.000 134.800 124.200 135.100 ;
        RECT 125.400 134.800 125.800 135.200 ;
        RECT 126.200 134.800 126.600 135.200 ;
        RECT 127.000 134.800 127.400 135.200 ;
        RECT 127.800 134.800 128.200 135.200 ;
        RECT 131.000 134.800 131.400 135.200 ;
        RECT 133.400 134.800 133.800 135.200 ;
        RECT 103.000 128.800 103.400 129.200 ;
        RECT 100.600 124.800 101.000 125.200 ;
        RECT 101.400 114.700 101.800 115.100 ;
        RECT 101.400 112.200 101.700 114.700 ;
        RECT 101.400 111.800 101.800 112.200 ;
        RECT 102.200 112.100 102.600 117.900 ;
        RECT 103.000 116.800 103.400 117.200 ;
        RECT 103.000 109.200 103.300 116.800 ;
        RECT 103.800 113.100 104.200 115.900 ;
        RECT 104.600 113.100 105.000 115.900 ;
        RECT 106.200 112.100 106.600 117.900 ;
        RECT 107.000 115.200 107.300 134.800 ;
        RECT 110.200 133.800 110.600 134.200 ;
        RECT 110.200 131.200 110.500 133.800 ;
        RECT 111.000 133.200 111.300 134.800 ;
        RECT 111.000 132.800 111.400 133.200 ;
        RECT 110.200 130.800 110.600 131.200 ;
        RECT 110.200 129.200 110.500 130.800 ;
        RECT 111.000 129.200 111.300 132.800 ;
        RECT 110.200 128.800 110.600 129.200 ;
        RECT 111.000 128.800 111.400 129.200 ;
        RECT 113.400 126.200 113.700 134.800 ;
        RECT 117.400 129.200 117.700 134.800 ;
        RECT 120.600 132.200 120.900 134.800 ;
        RECT 120.600 131.800 121.000 132.200 ;
        RECT 117.400 128.800 117.800 129.200 ;
        RECT 119.800 128.800 120.200 129.200 ;
        RECT 117.400 128.200 117.700 128.800 ;
        RECT 119.800 128.200 120.100 128.800 ;
        RECT 117.400 127.800 117.800 128.200 ;
        RECT 119.800 127.800 120.200 128.200 ;
        RECT 126.200 126.200 126.500 134.800 ;
        RECT 127.000 134.200 127.300 134.800 ;
        RECT 127.000 133.800 127.400 134.200 ;
        RECT 111.800 125.800 112.200 126.200 ;
        RECT 112.600 125.800 113.000 126.200 ;
        RECT 113.400 125.800 113.800 126.200 ;
        RECT 115.800 125.800 116.200 126.200 ;
        RECT 122.200 125.800 122.600 126.200 ;
        RECT 126.200 125.800 126.600 126.200 ;
        RECT 111.800 124.200 112.100 125.800 ;
        RECT 111.800 123.800 112.200 124.200 ;
        RECT 110.200 117.800 110.600 118.200 ;
        RECT 110.200 115.200 110.500 117.800 ;
        RECT 107.000 114.800 107.400 115.200 ;
        RECT 107.800 114.800 108.200 115.200 ;
        RECT 109.400 114.800 109.800 115.200 ;
        RECT 110.200 114.800 110.600 115.200 ;
        RECT 107.800 114.200 108.100 114.800 ;
        RECT 107.800 113.800 108.200 114.200 ;
        RECT 103.000 109.100 103.400 109.200 ;
        RECT 103.800 109.100 104.200 109.200 ;
        RECT 99.000 106.800 99.400 107.200 ;
        RECT 99.000 106.100 99.400 106.200 ;
        RECT 99.800 106.100 100.200 106.200 ;
        RECT 99.000 105.800 100.200 106.100 ;
        RECT 101.400 103.100 101.800 108.900 ;
        RECT 103.000 108.800 104.200 109.100 ;
        RECT 102.200 107.800 102.600 108.200 ;
        RECT 102.200 107.200 102.500 107.800 ;
        RECT 102.200 106.800 102.600 107.200 ;
        RECT 103.000 105.100 103.400 107.900 ;
        RECT 104.600 103.800 105.000 104.200 ;
        RECT 103.000 101.800 103.400 102.200 ;
        RECT 103.000 99.200 103.300 101.800 ;
        RECT 104.600 99.200 104.900 103.800 ;
        RECT 106.200 103.100 106.600 108.900 ;
        RECT 107.000 105.800 107.400 106.200 ;
        RECT 107.000 104.200 107.300 105.800 ;
        RECT 107.000 103.800 107.400 104.200 ;
        RECT 103.000 98.800 103.400 99.200 ;
        RECT 104.600 98.800 105.000 99.200 ;
        RECT 91.000 94.800 91.400 95.200 ;
        RECT 93.400 94.800 93.800 95.200 ;
        RECT 91.000 93.200 91.300 94.800 ;
        RECT 93.400 94.200 93.700 94.800 ;
        RECT 93.400 93.800 93.800 94.200 ;
        RECT 91.000 92.800 91.400 93.200 ;
        RECT 79.000 85.800 79.400 86.200 ;
        RECT 81.400 83.100 81.800 88.900 ;
        RECT 84.600 88.800 85.000 89.200 ;
        RECT 87.000 89.100 87.400 89.200 ;
        RECT 87.800 89.100 88.100 91.800 ;
        RECT 87.000 88.800 88.100 89.100 ;
        RECT 82.200 86.800 82.600 87.200 ;
        RECT 78.200 76.800 78.600 77.200 ;
        RECT 75.800 73.100 76.200 75.900 ;
        RECT 77.400 75.800 77.800 76.200 ;
        RECT 76.600 74.800 77.000 75.200 ;
        RECT 76.600 74.200 76.900 74.800 ;
        RECT 76.600 73.800 77.000 74.200 ;
        RECT 77.400 74.100 77.800 74.200 ;
        RECT 78.200 74.100 78.500 76.800 ;
        RECT 80.600 76.100 81.000 76.200 ;
        RECT 81.400 76.100 81.800 76.200 ;
        RECT 80.600 75.800 81.800 76.100 ;
        RECT 80.600 75.100 81.000 75.200 ;
        RECT 81.400 75.100 81.800 75.200 ;
        RECT 80.600 74.800 81.800 75.100 ;
        RECT 77.400 73.800 78.500 74.100 ;
        RECT 79.800 74.100 80.200 74.200 ;
        RECT 80.600 74.100 81.000 74.200 ;
        RECT 79.800 73.800 81.000 74.100 ;
        RECT 78.200 72.800 78.600 73.200 ;
        RECT 79.000 73.100 79.400 73.200 ;
        RECT 79.800 73.100 80.200 73.200 ;
        RECT 79.000 72.800 80.200 73.100 ;
        RECT 78.200 72.200 78.500 72.800 ;
        RECT 78.200 71.800 78.600 72.200 ;
        RECT 77.400 69.800 77.800 70.200 ;
        RECT 77.400 69.200 77.700 69.800 ;
        RECT 77.400 68.800 77.800 69.200 ;
        RECT 79.000 68.800 79.400 69.200 ;
        RECT 73.400 66.800 73.800 67.200 ;
        RECT 76.600 66.800 77.000 67.200 ;
        RECT 76.600 66.200 76.900 66.800 ;
        RECT 72.600 65.800 73.000 66.200 ;
        RECT 73.400 65.800 73.800 66.200 ;
        RECT 76.600 65.800 77.000 66.200 ;
        RECT 69.400 58.800 69.800 59.200 ;
        RECT 64.600 54.800 65.000 55.200 ;
        RECT 67.000 55.000 67.400 55.100 ;
        RECT 67.800 55.000 68.200 55.100 ;
        RECT 64.600 54.200 64.900 54.800 ;
        RECT 67.000 54.700 68.200 55.000 ;
        RECT 64.600 53.800 65.000 54.200 ;
        RECT 68.600 52.100 69.000 57.900 ;
        RECT 68.600 49.100 69.000 49.200 ;
        RECT 69.400 49.100 69.700 58.800 ;
        RECT 72.600 57.200 72.900 65.800 ;
        RECT 73.400 59.200 73.700 65.800 ;
        RECT 75.000 61.800 75.400 62.200 ;
        RECT 73.400 58.800 73.800 59.200 ;
        RECT 72.600 56.800 73.000 57.200 ;
        RECT 70.200 53.100 70.600 55.900 ;
        RECT 75.000 55.200 75.300 61.800 ;
        RECT 75.800 56.800 76.200 57.200 ;
        RECT 75.800 55.200 76.100 56.800 ;
        RECT 76.600 55.800 77.000 56.200 ;
        RECT 76.600 55.200 76.900 55.800 ;
        RECT 79.000 55.200 79.300 68.800 ;
        RECT 79.800 63.100 80.200 68.900 ;
        RECT 82.200 68.200 82.500 86.800 ;
        RECT 83.000 85.100 83.400 87.900 ;
        RECT 86.200 85.800 86.600 86.200 ;
        RECT 86.200 83.200 86.500 85.800 ;
        RECT 88.600 83.800 89.000 84.200 ;
        RECT 86.200 82.800 86.600 83.200 ;
        RECT 86.200 80.200 86.500 82.800 ;
        RECT 86.200 79.800 86.600 80.200 ;
        RECT 83.000 77.800 83.400 78.200 ;
        RECT 86.200 77.800 86.600 78.200 ;
        RECT 83.000 76.200 83.300 77.800 ;
        RECT 86.200 76.200 86.500 77.800 ;
        RECT 88.600 76.200 88.900 83.800 ;
        RECT 89.400 83.100 89.800 88.900 ;
        RECT 93.400 86.300 93.700 93.800 ;
        RECT 95.000 92.100 95.400 97.900 ;
        RECT 96.600 93.100 97.000 95.900 ;
        RECT 93.400 85.900 93.800 86.300 ;
        RECT 94.200 83.100 94.600 88.900 ;
        RECT 95.000 87.800 95.400 88.200 ;
        RECT 95.000 87.200 95.300 87.800 ;
        RECT 95.000 86.800 95.400 87.200 ;
        RECT 95.800 85.100 96.200 87.900 ;
        RECT 100.600 83.100 101.000 88.900 ;
        RECT 98.200 81.800 98.600 82.200 ;
        RECT 100.600 81.800 101.000 82.200 ;
        RECT 98.200 81.200 98.500 81.800 ;
        RECT 98.200 80.800 98.600 81.200 ;
        RECT 83.000 75.800 83.400 76.200 ;
        RECT 83.800 75.800 84.200 76.200 ;
        RECT 86.200 75.800 86.600 76.200 ;
        RECT 88.600 75.800 89.000 76.200 ;
        RECT 91.800 75.800 92.200 76.200 ;
        RECT 83.000 72.800 83.400 73.200 ;
        RECT 83.000 72.200 83.300 72.800 ;
        RECT 83.000 71.800 83.400 72.200 ;
        RECT 83.800 68.200 84.100 75.800 ;
        RECT 91.800 75.200 92.100 75.800 ;
        RECT 98.200 75.200 98.500 80.800 ;
        RECT 99.000 79.800 99.400 80.200 ;
        RECT 99.000 75.200 99.300 79.800 ;
        RECT 100.600 79.200 100.900 81.800 ;
        RECT 103.000 79.200 103.300 98.800 ;
        RECT 109.400 95.200 109.700 114.800 ;
        RECT 110.200 113.200 110.500 114.800 ;
        RECT 110.200 112.800 110.600 113.200 ;
        RECT 110.200 111.800 110.600 112.200 ;
        RECT 111.000 112.100 111.400 117.900 ;
        RECT 110.200 106.300 110.500 111.800 ;
        RECT 110.200 105.900 110.600 106.300 ;
        RECT 110.200 105.200 110.500 105.900 ;
        RECT 110.200 104.800 110.600 105.200 ;
        RECT 111.000 103.100 111.400 108.900 ;
        RECT 111.800 99.200 112.100 123.800 ;
        RECT 112.600 116.200 112.900 125.800 ;
        RECT 113.400 117.200 113.700 125.800 ;
        RECT 115.800 122.200 116.100 125.800 ;
        RECT 122.200 125.200 122.500 125.800 ;
        RECT 122.200 124.800 122.600 125.200 ;
        RECT 127.800 123.200 128.100 134.800 ;
        RECT 133.400 134.200 133.700 134.800 ;
        RECT 133.400 133.800 133.800 134.200 ;
        RECT 131.800 132.800 132.200 133.200 ;
        RECT 131.800 130.200 132.100 132.800 ;
        RECT 131.800 129.800 132.200 130.200 ;
        RECT 134.200 129.200 134.500 135.800 ;
        RECT 141.400 135.200 141.700 135.800 ;
        RECT 135.800 135.100 136.200 135.200 ;
        RECT 136.600 135.100 137.000 135.200 ;
        RECT 135.800 134.800 137.000 135.100 ;
        RECT 137.400 135.100 137.800 135.200 ;
        RECT 138.200 135.100 138.600 135.200 ;
        RECT 137.400 134.800 138.600 135.100 ;
        RECT 141.400 134.800 141.800 135.200 ;
        RECT 143.000 134.800 143.400 135.200 ;
        RECT 145.400 134.800 145.800 135.200 ;
        RECT 143.000 134.200 143.300 134.800 ;
        RECT 145.400 134.200 145.700 134.800 ;
        RECT 135.000 133.800 135.400 134.200 ;
        RECT 137.400 133.800 137.800 134.200 ;
        RECT 139.800 133.800 140.200 134.200 ;
        RECT 143.000 133.800 143.400 134.200 ;
        RECT 143.800 133.800 144.200 134.200 ;
        RECT 145.400 133.800 145.800 134.200 ;
        RECT 134.200 128.800 134.600 129.200 ;
        RECT 135.000 127.200 135.300 133.800 ;
        RECT 137.400 133.200 137.700 133.800 ;
        RECT 137.400 132.800 137.800 133.200 ;
        RECT 139.800 131.200 140.100 133.800 ;
        RECT 143.800 133.200 144.100 133.800 ;
        RECT 140.600 132.800 141.000 133.200 ;
        RECT 143.800 132.800 144.200 133.200 ;
        RECT 140.600 132.200 140.900 132.800 ;
        RECT 140.600 131.800 141.000 132.200 ;
        RECT 142.200 131.800 142.600 132.200 ;
        RECT 144.600 132.100 145.000 132.200 ;
        RECT 145.400 132.100 145.800 132.200 ;
        RECT 144.600 131.800 145.800 132.100 ;
        RECT 137.400 130.800 137.800 131.200 ;
        RECT 139.800 130.800 140.200 131.200 ;
        RECT 137.400 127.200 137.700 130.800 ;
        RECT 135.000 126.800 135.400 127.200 ;
        RECT 136.600 126.800 137.000 127.200 ;
        RECT 137.400 126.800 137.800 127.200 ;
        RECT 139.800 127.100 140.100 130.800 ;
        RECT 142.200 127.200 142.500 131.800 ;
        RECT 146.200 131.200 146.500 135.800 ;
        RECT 157.400 135.200 157.700 135.800 ;
        RECT 147.800 134.800 148.200 135.200 ;
        RECT 153.400 134.800 153.800 135.200 ;
        RECT 157.400 134.800 157.800 135.200 ;
        RECT 147.800 132.200 148.100 134.800 ;
        RECT 151.800 133.800 152.200 134.200 ;
        RECT 151.800 133.200 152.100 133.800 ;
        RECT 150.200 132.800 150.600 133.200 ;
        RECT 151.800 132.800 152.200 133.200 ;
        RECT 147.800 131.800 148.200 132.200 ;
        RECT 146.200 130.800 146.600 131.200 ;
        RECT 147.000 129.800 147.400 130.200 ;
        RECT 147.000 129.200 147.300 129.800 ;
        RECT 147.000 128.800 147.400 129.200 ;
        RECT 150.200 128.200 150.500 132.800 ;
        RECT 151.800 128.200 152.100 132.800 ;
        RECT 153.400 132.200 153.700 134.800 ;
        RECT 160.600 134.200 160.900 135.800 ;
        RECT 161.400 135.200 161.700 137.800 ;
        RECT 163.800 135.800 164.200 136.200 ;
        RECT 161.400 134.800 161.800 135.200 ;
        RECT 155.000 134.100 155.400 134.200 ;
        RECT 155.800 134.100 156.200 134.200 ;
        RECT 155.000 133.800 156.200 134.100 ;
        RECT 157.400 134.100 157.800 134.200 ;
        RECT 158.200 134.100 158.600 134.200 ;
        RECT 157.400 133.800 158.600 134.100 ;
        RECT 160.600 133.800 161.000 134.200 ;
        RECT 162.200 133.800 162.600 134.200 ;
        RECT 162.200 133.200 162.500 133.800 ;
        RECT 159.800 133.100 160.200 133.200 ;
        RECT 160.600 133.100 161.000 133.200 ;
        RECT 159.800 132.800 161.000 133.100 ;
        RECT 162.200 132.800 162.600 133.200 ;
        RECT 153.400 131.800 153.800 132.200 ;
        RECT 155.000 131.800 155.400 132.200 ;
        RECT 156.600 131.800 157.000 132.200 ;
        RECT 159.000 131.800 159.400 132.200 ;
        RECT 155.000 128.200 155.300 131.800 ;
        RECT 150.200 127.800 150.600 128.200 ;
        RECT 151.800 127.800 152.200 128.200 ;
        RECT 155.000 127.800 155.400 128.200 ;
        RECT 139.800 126.800 140.900 127.100 ;
        RECT 142.200 126.800 142.600 127.200 ;
        RECT 143.000 126.800 143.400 127.200 ;
        RECT 143.800 126.800 144.200 127.200 ;
        RECT 129.400 125.800 129.800 126.200 ;
        RECT 132.600 125.800 133.000 126.200 ;
        RECT 129.400 125.200 129.700 125.800 ;
        RECT 129.400 124.800 129.800 125.200 ;
        RECT 132.600 124.200 132.900 125.800 ;
        RECT 132.600 123.800 133.000 124.200 ;
        RECT 127.800 122.800 128.200 123.200 ;
        RECT 115.000 121.800 115.400 122.200 ;
        RECT 115.800 121.800 116.200 122.200 ;
        RECT 126.200 121.800 126.600 122.200 ;
        RECT 127.800 121.800 128.200 122.200 ;
        RECT 131.000 121.800 131.400 122.200 ;
        RECT 113.400 116.800 113.800 117.200 ;
        RECT 114.200 116.800 114.600 117.200 ;
        RECT 112.600 115.800 113.000 116.200 ;
        RECT 112.600 111.200 112.900 115.800 ;
        RECT 114.200 115.200 114.500 116.800 ;
        RECT 114.200 114.800 114.600 115.200 ;
        RECT 113.400 112.800 113.800 113.200 ;
        RECT 112.600 110.800 113.000 111.200 ;
        RECT 113.400 108.200 113.700 112.800 ;
        RECT 112.600 105.100 113.000 107.900 ;
        RECT 113.400 107.800 113.800 108.200 ;
        RECT 113.400 106.800 113.800 107.200 ;
        RECT 113.400 106.200 113.700 106.800 ;
        RECT 115.000 106.200 115.300 121.800 ;
        RECT 116.600 112.100 117.000 117.900 ;
        RECT 117.400 114.800 117.800 115.200 ;
        RECT 117.400 111.100 117.700 114.800 ;
        RECT 120.600 114.700 121.000 115.100 ;
        RECT 120.600 114.200 120.900 114.700 ;
        RECT 120.600 113.800 121.000 114.200 ;
        RECT 121.400 112.100 121.800 117.900 ;
        RECT 123.800 117.800 124.200 118.200 ;
        RECT 123.000 113.100 123.400 115.900 ;
        RECT 123.800 113.200 124.100 117.800 ;
        RECT 125.400 115.800 125.800 116.200 ;
        RECT 125.400 115.200 125.700 115.800 ;
        RECT 126.200 115.200 126.500 121.800 ;
        RECT 127.800 118.200 128.100 121.800 ;
        RECT 131.000 118.200 131.300 121.800 ;
        RECT 127.800 118.100 128.200 118.200 ;
        RECT 127.800 117.800 128.900 118.100 ;
        RECT 131.000 117.800 131.400 118.200 ;
        RECT 127.800 116.800 128.200 117.200 ;
        RECT 127.800 116.200 128.100 116.800 ;
        RECT 127.800 115.800 128.200 116.200 ;
        RECT 125.400 114.800 125.800 115.200 ;
        RECT 126.200 114.800 126.600 115.200 ;
        RECT 124.600 114.100 125.000 114.200 ;
        RECT 125.400 114.100 125.800 114.200 ;
        RECT 124.600 113.800 125.800 114.100 ;
        RECT 123.800 112.800 124.200 113.200 ;
        RECT 123.800 111.800 124.200 112.200 ;
        RECT 116.600 110.800 117.700 111.100 ;
        RECT 123.000 110.800 123.400 111.200 ;
        RECT 116.600 109.200 116.900 110.800 ;
        RECT 121.400 109.800 121.800 110.200 ;
        RECT 116.600 108.800 117.000 109.200 ;
        RECT 116.600 107.200 116.900 108.800 ;
        RECT 116.600 106.800 117.000 107.200 ;
        RECT 113.400 105.800 113.800 106.200 ;
        RECT 115.000 105.800 115.400 106.200 ;
        RECT 111.800 98.800 112.200 99.200 ;
        RECT 118.200 98.800 118.600 99.200 ;
        RECT 111.800 97.800 112.200 98.200 ;
        RECT 115.800 97.800 116.200 98.200 ;
        RECT 111.800 95.200 112.100 97.800 ;
        RECT 113.400 95.800 113.800 96.200 ;
        RECT 107.800 94.800 108.200 95.200 ;
        RECT 108.600 94.800 109.000 95.200 ;
        RECT 109.400 94.800 109.800 95.200 ;
        RECT 111.800 94.800 112.200 95.200 ;
        RECT 107.800 94.200 108.100 94.800 ;
        RECT 107.800 93.800 108.200 94.200 ;
        RECT 105.400 93.100 105.800 93.200 ;
        RECT 106.200 93.100 106.600 93.200 ;
        RECT 105.400 92.800 106.600 93.100 ;
        RECT 104.600 91.800 105.000 92.200 ;
        RECT 107.000 91.800 107.400 92.200 ;
        RECT 104.600 87.200 104.900 91.800 ;
        RECT 107.000 89.200 107.300 91.800 ;
        RECT 104.600 86.800 105.000 87.200 ;
        RECT 104.600 85.900 105.000 86.300 ;
        RECT 104.600 85.200 104.900 85.900 ;
        RECT 104.600 84.800 105.000 85.200 ;
        RECT 105.400 83.100 105.800 88.900 ;
        RECT 107.000 88.800 107.400 89.200 ;
        RECT 106.200 87.800 106.600 88.200 ;
        RECT 106.200 87.200 106.500 87.800 ;
        RECT 106.200 86.800 106.600 87.200 ;
        RECT 99.800 78.800 100.200 79.200 ;
        RECT 100.600 78.800 101.000 79.200 ;
        RECT 103.000 78.800 103.400 79.200 ;
        RECT 84.600 75.100 85.000 75.200 ;
        RECT 85.400 75.100 85.800 75.200 ;
        RECT 84.600 74.800 85.800 75.100 ;
        RECT 87.800 74.800 88.200 75.200 ;
        RECT 88.600 74.800 89.000 75.200 ;
        RECT 91.800 74.800 92.200 75.200 ;
        RECT 92.600 75.100 93.000 75.200 ;
        RECT 93.400 75.100 93.800 75.200 ;
        RECT 92.600 74.800 93.800 75.100 ;
        RECT 95.800 74.800 96.200 75.200 ;
        RECT 96.600 74.800 97.000 75.200 ;
        RECT 98.200 74.800 98.600 75.200 ;
        RECT 99.000 74.800 99.400 75.200 ;
        RECT 85.400 74.100 85.800 74.200 ;
        RECT 86.200 74.100 86.600 74.200 ;
        RECT 85.400 73.800 86.600 74.100 ;
        RECT 86.200 71.800 86.600 72.200 ;
        RECT 86.200 71.200 86.500 71.800 ;
        RECT 86.200 70.800 86.600 71.200 ;
        RECT 87.800 69.200 88.100 74.800 ;
        RECT 88.600 74.200 88.900 74.800 ;
        RECT 88.600 73.800 89.000 74.200 ;
        RECT 94.200 71.800 94.600 72.200 ;
        RECT 94.200 69.200 94.500 71.800 ;
        RECT 95.800 70.200 96.100 74.800 ;
        RECT 96.600 72.200 96.900 74.800 ;
        RECT 96.600 71.800 97.000 72.200 ;
        RECT 95.800 69.800 96.200 70.200 ;
        RECT 99.800 69.200 100.100 78.800 ;
        RECT 103.000 76.200 103.300 78.800 ;
        RECT 106.200 77.100 106.500 86.800 ;
        RECT 107.000 85.100 107.400 87.900 ;
        RECT 108.600 86.200 108.900 94.800 ;
        RECT 109.400 88.200 109.700 94.800 ;
        RECT 113.400 94.200 113.700 95.800 ;
        RECT 115.000 94.800 115.400 95.200 ;
        RECT 110.200 93.800 110.600 94.200 ;
        RECT 113.400 93.800 113.800 94.200 ;
        RECT 110.200 93.200 110.500 93.800 ;
        RECT 110.200 92.800 110.600 93.200 ;
        RECT 115.000 92.200 115.300 94.800 ;
        RECT 115.800 94.200 116.100 97.800 ;
        RECT 118.200 94.200 118.500 98.800 ;
        RECT 119.000 98.100 119.400 98.200 ;
        RECT 119.800 98.100 120.200 98.200 ;
        RECT 119.000 97.800 120.200 98.100 ;
        RECT 120.600 95.800 121.000 96.200 ;
        RECT 115.800 93.800 116.200 94.200 ;
        RECT 116.600 94.100 117.000 94.200 ;
        RECT 117.400 94.100 117.800 94.200 ;
        RECT 116.600 93.800 117.800 94.100 ;
        RECT 118.200 93.800 118.600 94.200 ;
        RECT 119.800 93.800 120.200 94.200 ;
        RECT 119.800 93.200 120.100 93.800 ;
        RECT 119.800 92.800 120.200 93.200 ;
        RECT 115.000 91.800 115.400 92.200 ;
        RECT 119.800 91.800 120.200 92.200 ;
        RECT 109.400 87.800 109.800 88.200 ;
        RECT 108.600 85.800 109.000 86.200 ;
        RECT 107.800 81.800 108.200 82.200 ;
        RECT 107.800 81.200 108.100 81.800 ;
        RECT 107.800 80.800 108.200 81.200 ;
        RECT 106.200 76.800 107.300 77.100 ;
        RECT 103.000 75.800 103.400 76.200 ;
        RECT 105.400 73.800 105.800 74.200 ;
        RECT 82.200 67.800 82.600 68.200 ;
        RECT 83.800 67.800 84.200 68.200 ;
        RECT 83.000 66.200 83.400 66.300 ;
        RECT 83.800 66.200 84.200 66.300 ;
        RECT 83.000 65.900 84.200 66.200 ;
        RECT 84.600 63.100 85.000 68.900 ;
        RECT 87.800 68.800 88.200 69.200 ;
        RECT 88.600 68.800 89.000 69.200 ;
        RECT 87.000 68.100 87.400 68.200 ;
        RECT 87.800 68.100 88.200 68.200 ;
        RECT 86.200 65.100 86.600 67.900 ;
        RECT 87.000 67.800 88.200 68.100 ;
        RECT 88.600 66.200 88.900 68.800 ;
        RECT 87.000 66.100 87.400 66.200 ;
        RECT 87.800 66.100 88.200 66.200 ;
        RECT 87.000 65.800 88.200 66.100 ;
        RECT 88.600 65.800 89.000 66.200 ;
        RECT 89.400 65.100 89.800 67.900 ;
        RECT 91.000 63.100 91.400 68.900 ;
        RECT 94.200 68.800 94.600 69.200 ;
        RECT 97.400 69.100 97.800 69.200 ;
        RECT 98.200 69.100 98.600 69.200 ;
        RECT 93.400 67.800 93.800 68.200 ;
        RECT 93.400 67.200 93.700 67.800 ;
        RECT 91.800 66.800 92.200 67.200 ;
        RECT 93.400 67.100 93.800 67.200 ;
        RECT 94.200 67.100 94.600 67.200 ;
        RECT 93.400 66.800 94.600 67.100 ;
        RECT 91.800 66.300 92.100 66.800 ;
        RECT 91.800 65.900 92.200 66.300 ;
        RECT 95.800 63.100 96.200 68.900 ;
        RECT 97.400 68.800 98.600 69.100 ;
        RECT 99.800 68.800 100.200 69.200 ;
        RECT 103.000 63.100 103.400 68.900 ;
        RECT 103.800 67.800 104.200 68.200 ;
        RECT 103.800 67.200 104.100 67.800 ;
        RECT 103.800 66.800 104.200 67.200 ;
        RECT 105.400 57.200 105.700 73.800 ;
        RECT 106.200 73.100 106.600 75.900 ;
        RECT 107.000 68.200 107.300 76.800 ;
        RECT 107.800 72.100 108.200 77.900 ;
        RECT 108.600 72.200 108.900 85.800 ;
        RECT 110.200 83.100 110.600 88.900 ;
        RECT 113.400 88.800 113.800 89.200 ;
        RECT 114.200 88.800 114.600 89.200 ;
        RECT 111.000 86.800 111.400 87.200 ;
        RECT 111.000 86.200 111.300 86.800 ;
        RECT 113.400 86.200 113.700 88.800 ;
        RECT 111.000 85.800 111.400 86.200 ;
        RECT 113.400 85.800 113.800 86.200 ;
        RECT 111.000 75.200 111.300 85.800 ;
        RECT 114.200 79.200 114.500 88.800 ;
        RECT 115.000 83.100 115.400 88.900 ;
        RECT 116.600 85.100 117.000 87.900 ;
        RECT 117.400 87.800 117.800 88.200 ;
        RECT 117.400 79.200 117.700 87.800 ;
        RECT 119.000 86.800 119.400 87.200 ;
        RECT 119.000 86.200 119.300 86.800 ;
        RECT 119.000 85.800 119.400 86.200 ;
        RECT 119.800 85.200 120.100 91.800 ;
        RECT 120.600 89.200 120.900 95.800 ;
        RECT 121.400 95.200 121.700 109.800 ;
        RECT 123.000 106.200 123.300 110.800 ;
        RECT 123.800 106.200 124.100 111.800 ;
        RECT 126.200 110.800 126.600 111.200 ;
        RECT 124.600 108.800 125.000 109.200 ;
        RECT 123.000 105.800 123.400 106.200 ;
        RECT 123.800 105.800 124.200 106.200 ;
        RECT 121.400 95.100 121.800 95.200 ;
        RECT 122.200 95.100 122.600 95.200 ;
        RECT 121.400 94.800 122.600 95.100 ;
        RECT 123.000 94.100 123.300 105.800 ;
        RECT 122.200 93.800 123.300 94.100 ;
        RECT 120.600 88.800 121.000 89.200 ;
        RECT 121.400 87.800 121.800 88.200 ;
        RECT 121.400 87.200 121.700 87.800 ;
        RECT 121.400 86.800 121.800 87.200 ;
        RECT 122.200 86.200 122.500 93.800 ;
        RECT 123.800 89.200 124.100 105.800 ;
        RECT 124.600 93.200 124.900 108.800 ;
        RECT 126.200 106.200 126.500 110.800 ;
        RECT 126.200 105.800 126.600 106.200 ;
        RECT 127.800 105.100 128.200 107.900 ;
        RECT 128.600 107.200 128.900 117.800 ;
        RECT 131.000 116.800 131.400 117.200 ;
        RECT 131.000 116.200 131.300 116.800 ;
        RECT 131.000 115.800 131.400 116.200 ;
        RECT 135.000 115.200 135.300 126.800 ;
        RECT 136.600 126.200 136.900 126.800 ;
        RECT 136.600 125.800 137.000 126.200 ;
        RECT 138.200 125.800 138.600 126.200 ;
        RECT 138.200 125.200 138.500 125.800 ;
        RECT 138.200 124.800 138.600 125.200 ;
        RECT 139.000 125.100 139.400 125.200 ;
        RECT 139.800 125.100 140.200 125.200 ;
        RECT 139.000 124.800 140.200 125.100 ;
        RECT 140.600 121.200 140.900 126.800 ;
        RECT 143.000 126.200 143.300 126.800 ;
        RECT 143.800 126.200 144.100 126.800 ;
        RECT 150.200 126.200 150.500 127.800 ;
        RECT 141.400 125.800 141.800 126.200 ;
        RECT 143.000 125.800 143.400 126.200 ;
        RECT 143.800 125.800 144.200 126.200 ;
        RECT 145.400 126.100 145.800 126.200 ;
        RECT 146.200 126.100 146.600 126.200 ;
        RECT 145.400 125.800 146.600 126.100 ;
        RECT 147.800 125.800 148.200 126.200 ;
        RECT 150.200 125.800 150.600 126.200 ;
        RECT 140.600 120.800 141.000 121.200 ;
        RECT 135.800 115.800 136.200 116.200 ;
        RECT 137.400 115.800 137.800 116.200 ;
        RECT 129.400 114.800 129.800 115.200 ;
        RECT 130.200 115.100 130.600 115.200 ;
        RECT 131.000 115.100 131.400 115.200 ;
        RECT 130.200 114.800 131.400 115.100 ;
        RECT 135.000 114.800 135.400 115.200 ;
        RECT 129.400 114.200 129.700 114.800 ;
        RECT 135.800 114.200 136.100 115.800 ;
        RECT 137.400 115.200 137.700 115.800 ;
        RECT 137.400 114.800 137.800 115.200 ;
        RECT 139.800 114.800 140.200 115.200 ;
        RECT 129.400 113.800 129.800 114.200 ;
        RECT 135.000 114.100 135.400 114.200 ;
        RECT 135.800 114.100 136.200 114.200 ;
        RECT 135.000 113.800 136.200 114.100 ;
        RECT 133.400 112.800 133.800 113.200 ;
        RECT 131.800 111.800 132.200 112.200 ;
        RECT 128.600 106.800 129.000 107.200 ;
        RECT 129.400 103.100 129.800 108.900 ;
        RECT 130.200 106.100 130.600 106.200 ;
        RECT 131.000 106.100 131.400 106.200 ;
        RECT 130.200 105.800 131.400 106.100 ;
        RECT 125.400 101.800 125.800 102.200 ;
        RECT 125.400 95.200 125.700 101.800 ;
        RECT 131.800 97.200 132.100 111.800 ;
        RECT 133.400 109.200 133.700 112.800 ;
        RECT 137.400 110.200 137.700 114.800 ;
        RECT 139.800 114.200 140.100 114.800 ;
        RECT 139.800 113.800 140.200 114.200 ;
        RECT 137.400 109.800 137.800 110.200 ;
        RECT 133.400 108.800 133.800 109.200 ;
        RECT 135.800 109.100 136.200 109.200 ;
        RECT 136.600 109.100 137.000 109.200 ;
        RECT 134.200 103.100 134.600 108.900 ;
        RECT 135.800 108.800 137.000 109.100 ;
        RECT 135.000 106.800 135.400 107.200 ;
        RECT 131.800 96.800 132.200 97.200 ;
        RECT 133.400 96.800 133.800 97.200 ;
        RECT 126.200 95.900 126.600 96.300 ;
        RECT 129.300 95.900 129.700 96.300 ;
        RECT 125.400 94.800 125.800 95.200 ;
        RECT 126.200 94.200 126.500 95.900 ;
        RECT 128.700 94.900 129.100 95.300 ;
        RECT 128.700 94.200 129.000 94.900 ;
        RECT 125.400 93.800 125.800 94.200 ;
        RECT 126.200 93.900 129.000 94.200 ;
        RECT 125.400 93.200 125.700 93.800 ;
        RECT 126.200 93.500 126.500 93.900 ;
        RECT 126.900 93.500 127.300 93.600 ;
        RECT 128.600 93.500 129.000 93.600 ;
        RECT 129.400 93.500 129.700 95.900 ;
        RECT 133.400 95.200 133.700 96.800 ;
        RECT 133.400 94.800 133.800 95.200 ;
        RECT 130.200 94.100 130.600 94.200 ;
        RECT 131.000 94.100 131.400 94.200 ;
        RECT 130.200 93.800 131.400 94.100 ;
        RECT 133.400 93.800 133.800 94.200 ;
        RECT 124.600 92.800 125.000 93.200 ;
        RECT 125.400 92.800 125.800 93.200 ;
        RECT 126.200 93.100 126.600 93.500 ;
        RECT 126.900 93.200 129.700 93.500 ;
        RECT 129.300 93.100 129.700 93.200 ;
        RECT 131.000 92.800 131.400 93.200 ;
        RECT 131.000 92.200 131.300 92.800 ;
        RECT 133.400 92.200 133.700 93.800 ;
        RECT 127.800 92.100 128.200 92.200 ;
        RECT 128.600 92.100 129.000 92.200 ;
        RECT 127.800 91.800 129.000 92.100 ;
        RECT 131.000 91.800 131.400 92.200 ;
        RECT 131.800 92.100 132.200 92.200 ;
        RECT 132.600 92.100 133.000 92.200 ;
        RECT 131.800 91.800 133.000 92.100 ;
        RECT 133.400 91.800 133.800 92.200 ;
        RECT 123.800 88.800 124.200 89.200 ;
        RECT 127.000 88.800 127.400 89.200 ;
        RECT 127.000 88.200 127.300 88.800 ;
        RECT 123.800 87.800 124.200 88.200 ;
        RECT 127.000 87.800 127.400 88.200 ;
        RECT 123.800 87.200 124.100 87.800 ;
        RECT 123.800 86.800 124.200 87.200 ;
        RECT 121.400 86.100 121.800 86.200 ;
        RECT 122.200 86.100 122.600 86.200 ;
        RECT 121.400 85.800 122.600 86.100 ;
        RECT 123.000 85.800 123.400 86.200 ;
        RECT 125.400 86.100 125.800 86.200 ;
        RECT 126.200 86.100 126.600 86.200 ;
        RECT 125.400 85.800 126.600 86.100 ;
        RECT 119.800 84.800 120.200 85.200 ;
        RECT 119.800 82.200 120.100 84.800 ;
        RECT 119.000 81.800 119.400 82.200 ;
        RECT 119.800 81.800 120.200 82.200 ;
        RECT 114.200 79.100 114.600 79.200 ;
        RECT 115.000 79.100 115.400 79.200 ;
        RECT 114.200 78.800 115.400 79.100 ;
        RECT 117.400 78.800 117.800 79.200 ;
        RECT 109.400 74.800 109.800 75.200 ;
        RECT 111.000 74.800 111.400 75.200 ;
        RECT 109.400 73.200 109.700 74.800 ;
        RECT 111.000 74.200 111.300 74.800 ;
        RECT 111.000 73.800 111.400 74.200 ;
        RECT 109.400 72.800 109.800 73.200 ;
        RECT 108.600 71.800 109.000 72.200 ;
        RECT 111.000 71.800 111.400 72.200 ;
        RECT 112.600 72.100 113.000 77.900 ;
        RECT 115.800 73.100 116.200 75.900 ;
        RECT 116.600 73.800 117.000 74.200 ;
        RECT 107.000 67.800 107.400 68.200 ;
        RECT 107.000 66.800 107.400 67.200 ;
        RECT 107.000 66.300 107.300 66.800 ;
        RECT 107.000 65.900 107.400 66.300 ;
        RECT 107.800 63.100 108.200 68.900 ;
        RECT 109.400 65.100 109.800 67.900 ;
        RECT 111.000 59.200 111.300 71.800 ;
        RECT 116.600 69.200 116.900 73.800 ;
        RECT 117.400 72.100 117.800 77.900 ;
        RECT 119.000 75.200 119.300 81.800 ;
        RECT 121.400 78.800 121.800 79.200 ;
        RECT 121.400 76.200 121.700 78.800 ;
        RECT 121.400 75.800 121.800 76.200 ;
        RECT 121.400 75.200 121.700 75.800 ;
        RECT 119.000 74.800 119.400 75.200 ;
        RECT 121.400 74.800 121.800 75.200 ;
        RECT 113.400 67.800 113.800 68.200 ;
        RECT 113.400 66.200 113.700 67.800 ;
        RECT 113.400 65.800 113.800 66.200 ;
        RECT 114.200 65.100 114.600 67.900 ;
        RECT 115.800 63.100 116.200 68.900 ;
        RECT 116.600 68.800 117.000 69.200 ;
        RECT 116.600 68.200 116.900 68.800 ;
        RECT 116.600 67.800 117.000 68.200 ;
        RECT 119.000 66.200 119.300 74.800 ;
        RECT 122.200 72.100 122.600 77.900 ;
        RECT 123.000 76.200 123.300 85.800 ;
        RECT 129.400 83.100 129.800 88.900 ;
        RECT 132.600 86.800 133.000 87.200 ;
        RECT 133.400 86.800 133.800 87.200 ;
        RECT 132.600 86.200 132.900 86.800 ;
        RECT 132.600 85.800 133.000 86.200 ;
        RECT 123.000 75.800 123.400 76.200 ;
        RECT 127.000 75.800 127.400 76.200 ;
        RECT 125.400 75.100 125.800 75.200 ;
        RECT 126.200 75.100 126.600 75.200 ;
        RECT 125.400 74.800 126.600 75.100 ;
        RECT 125.400 73.800 125.800 74.200 ;
        RECT 125.400 73.200 125.700 73.800 ;
        RECT 127.000 73.200 127.300 75.800 ;
        RECT 125.400 72.800 125.800 73.200 ;
        RECT 127.000 73.100 127.400 73.200 ;
        RECT 127.800 73.100 128.200 73.200 ;
        RECT 127.000 72.800 128.200 73.100 ;
        RECT 124.600 71.800 125.000 72.200 ;
        RECT 119.000 65.800 119.400 66.200 ;
        RECT 120.600 63.100 121.000 68.900 ;
        RECT 124.600 64.200 124.900 71.800 ;
        RECT 133.400 69.200 133.700 86.800 ;
        RECT 134.200 83.100 134.600 88.900 ;
        RECT 135.000 87.200 135.300 106.800 ;
        RECT 137.400 105.100 137.800 107.900 ;
        RECT 138.200 107.800 138.600 108.200 ;
        RECT 138.200 107.200 138.500 107.800 ;
        RECT 138.200 106.800 138.600 107.200 ;
        RECT 139.000 103.100 139.400 108.900 ;
        RECT 141.400 106.200 141.700 125.800 ;
        RECT 143.000 120.800 143.400 121.200 ;
        RECT 143.000 119.200 143.300 120.800 ;
        RECT 143.000 118.800 143.400 119.200 ;
        RECT 142.200 114.800 142.600 115.200 ;
        RECT 142.200 113.200 142.500 114.800 ;
        RECT 142.200 112.800 142.600 113.200 ;
        RECT 143.800 111.100 144.100 125.800 ;
        RECT 147.800 125.200 148.100 125.800 ;
        RECT 145.400 124.800 145.800 125.200 ;
        RECT 147.800 124.800 148.200 125.200 ;
        RECT 145.400 121.200 145.700 124.800 ;
        RECT 150.200 121.800 150.600 122.200 ;
        RECT 145.400 120.800 145.800 121.200 ;
        RECT 143.000 110.800 144.100 111.100 ;
        RECT 145.400 112.800 145.800 113.200 ;
        RECT 142.200 108.800 142.600 109.200 ;
        RECT 141.400 105.800 141.800 106.200 ;
        RECT 138.300 95.900 138.700 96.300 ;
        RECT 141.400 95.900 141.800 96.300 ;
        RECT 137.400 93.800 137.800 94.200 ;
        RECT 137.400 88.200 137.700 93.800 ;
        RECT 138.300 93.500 138.600 95.900 ;
        RECT 138.900 94.900 139.300 95.300 ;
        RECT 139.000 94.200 139.300 94.900 ;
        RECT 141.500 94.200 141.800 95.900 ;
        RECT 139.000 93.900 141.800 94.200 ;
        RECT 139.000 93.500 139.400 93.600 ;
        RECT 140.700 93.500 141.100 93.600 ;
        RECT 141.500 93.500 141.800 93.900 ;
        RECT 142.200 94.200 142.500 108.800 ;
        RECT 143.000 99.200 143.300 110.800 ;
        RECT 145.400 109.200 145.700 112.800 ;
        RECT 146.200 111.800 146.600 112.200 ;
        RECT 148.600 112.100 149.000 117.900 ;
        RECT 150.200 117.200 150.500 121.800 ;
        RECT 150.200 116.800 150.600 117.200 ;
        RECT 151.800 115.200 152.100 127.800 ;
        RECT 152.600 126.800 153.000 127.200 ;
        RECT 155.000 126.800 155.400 127.200 ;
        RECT 152.600 126.200 152.900 126.800 ;
        RECT 155.000 126.200 155.300 126.800 ;
        RECT 152.600 125.800 153.000 126.200 ;
        RECT 155.000 125.800 155.400 126.200 ;
        RECT 155.800 124.800 156.200 125.200 ;
        RECT 155.800 124.200 156.100 124.800 ;
        RECT 156.600 124.200 156.900 131.800 ;
        RECT 159.000 129.100 159.300 131.800 ;
        RECT 159.000 128.800 160.100 129.100 ;
        RECT 159.000 127.800 159.400 128.200 ;
        RECT 159.000 127.200 159.300 127.800 ;
        RECT 157.400 126.800 157.800 127.200 ;
        RECT 159.000 126.800 159.400 127.200 ;
        RECT 157.400 126.200 157.700 126.800 ;
        RECT 157.400 125.800 157.800 126.200 ;
        RECT 157.400 124.200 157.700 125.800 ;
        RECT 158.200 125.100 158.600 125.200 ;
        RECT 159.000 125.100 159.400 125.200 ;
        RECT 158.200 124.800 159.400 125.100 ;
        RECT 155.800 123.800 156.200 124.200 ;
        RECT 156.600 123.800 157.000 124.200 ;
        RECT 157.400 123.800 157.800 124.200 ;
        RECT 151.800 114.800 152.200 115.200 ;
        RECT 152.600 114.700 153.000 115.100 ;
        RECT 149.400 113.800 149.800 114.200 ;
        RECT 146.200 110.200 146.500 111.800 ;
        RECT 146.200 109.800 146.600 110.200 ;
        RECT 147.000 109.800 147.400 110.200 ;
        RECT 145.400 109.100 145.800 109.200 ;
        RECT 146.200 109.100 146.600 109.200 ;
        RECT 143.800 103.100 144.200 108.900 ;
        RECT 145.400 108.800 146.600 109.100 ;
        RECT 147.000 107.200 147.300 109.800 ;
        RECT 147.000 106.800 147.400 107.200 ;
        RECT 149.400 106.200 149.700 113.800 ;
        RECT 152.600 112.200 152.900 114.700 ;
        RECT 152.600 111.800 153.000 112.200 ;
        RECT 153.400 112.100 153.800 117.900 ;
        RECT 154.200 113.800 154.600 114.200 ;
        RECT 154.200 113.200 154.500 113.800 ;
        RECT 154.200 112.800 154.600 113.200 ;
        RECT 155.000 113.100 155.400 115.900 ;
        RECT 155.800 115.800 156.200 116.200 ;
        RECT 156.600 115.800 157.000 116.200 ;
        RECT 155.800 114.200 156.100 115.800 ;
        RECT 156.600 115.200 156.900 115.800 ;
        RECT 156.600 115.100 157.000 115.200 ;
        RECT 156.600 114.800 157.700 115.100 ;
        RECT 155.800 113.800 156.200 114.200 ;
        RECT 152.600 106.800 153.000 107.200 ;
        RECT 152.600 106.200 152.900 106.800 ;
        RECT 149.400 105.800 149.800 106.200 ;
        RECT 152.600 105.800 153.000 106.200 ;
        RECT 149.400 105.200 149.700 105.800 ;
        RECT 149.400 104.800 149.800 105.200 ;
        RECT 154.200 102.200 154.500 112.800 ;
        RECT 155.000 108.800 155.400 109.200 ;
        RECT 155.000 108.200 155.300 108.800 ;
        RECT 155.800 108.200 156.100 113.800 ;
        RECT 155.000 107.800 155.400 108.200 ;
        RECT 155.800 107.800 156.200 108.200 ;
        RECT 157.400 106.200 157.700 114.800 ;
        RECT 158.200 111.800 158.600 112.200 ;
        RECT 159.000 111.800 159.400 112.200 ;
        RECT 158.200 107.200 158.500 111.800 ;
        RECT 159.000 110.200 159.300 111.800 ;
        RECT 159.000 109.800 159.400 110.200 ;
        RECT 158.200 106.800 158.600 107.200 ;
        RECT 155.800 106.100 156.200 106.200 ;
        RECT 156.600 106.100 157.000 106.200 ;
        RECT 155.800 105.800 157.000 106.100 ;
        RECT 157.400 105.800 157.800 106.200 ;
        RECT 158.200 106.100 158.600 106.200 ;
        RECT 159.000 106.100 159.400 106.200 ;
        RECT 158.200 105.800 159.400 106.100 ;
        RECT 151.000 101.800 151.400 102.200 ;
        RECT 154.200 101.800 154.600 102.200 ;
        RECT 159.000 101.800 159.400 102.200 ;
        RECT 143.000 98.800 143.400 99.200 ;
        RECT 142.200 93.800 142.600 94.200 ;
        RECT 143.000 93.800 143.400 94.200 ;
        RECT 138.300 93.200 141.100 93.500 ;
        RECT 138.300 93.100 138.700 93.200 ;
        RECT 141.400 93.100 141.800 93.500 ;
        RECT 143.000 93.200 143.300 93.800 ;
        RECT 143.000 92.800 143.400 93.200 ;
        RECT 139.000 92.100 139.400 92.200 ;
        RECT 139.800 92.100 140.200 92.200 ;
        RECT 145.400 92.100 145.800 97.900 ;
        RECT 149.400 95.800 149.800 96.200 ;
        RECT 149.400 95.100 149.700 95.800 ;
        RECT 149.400 94.700 149.800 95.100 ;
        RECT 150.200 92.100 150.600 97.900 ;
        RECT 151.000 94.200 151.300 101.800 ;
        RECT 153.400 99.100 153.800 99.200 ;
        RECT 154.200 99.100 154.600 99.200 ;
        RECT 153.400 98.800 154.600 99.100 ;
        RECT 151.000 93.800 151.400 94.200 ;
        RECT 139.000 91.800 140.200 92.100 ;
        RECT 143.000 90.800 143.400 91.200 ;
        RECT 135.000 86.800 135.400 87.200 ;
        RECT 135.800 85.100 136.200 87.900 ;
        RECT 136.600 87.800 137.000 88.200 ;
        RECT 137.400 87.800 137.800 88.200 ;
        RECT 142.200 87.800 142.600 88.200 ;
        RECT 136.600 74.200 136.900 87.800 ;
        RECT 137.400 87.100 137.800 87.200 ;
        RECT 138.200 87.100 138.600 87.200 ;
        RECT 137.400 86.800 138.600 87.100 ;
        RECT 139.000 86.800 139.400 87.200 ;
        RECT 139.000 86.200 139.300 86.800 ;
        RECT 142.200 86.200 142.500 87.800 ;
        RECT 143.000 86.200 143.300 90.800 ;
        RECT 145.400 88.800 145.800 89.200 ;
        RECT 145.400 88.200 145.700 88.800 ;
        RECT 145.400 87.800 145.800 88.200 ;
        RECT 138.200 85.800 138.600 86.200 ;
        RECT 139.000 85.800 139.400 86.200 ;
        RECT 140.600 85.800 141.000 86.200 ;
        RECT 142.200 85.800 142.600 86.200 ;
        RECT 143.000 85.800 143.400 86.200 ;
        RECT 138.200 85.200 138.500 85.800 ;
        RECT 140.600 85.200 140.900 85.800 ;
        RECT 138.200 84.800 138.600 85.200 ;
        RECT 140.600 84.800 141.000 85.200 ;
        RECT 137.400 83.800 137.800 84.200 ;
        RECT 137.400 79.200 137.700 83.800 ;
        RECT 147.800 83.100 148.200 88.900 ;
        RECT 151.000 87.200 151.300 93.800 ;
        RECT 151.800 93.100 152.200 95.900 ;
        RECT 156.600 92.100 157.000 97.900 ;
        RECT 159.000 97.200 159.300 101.800 ;
        RECT 159.000 96.800 159.400 97.200 ;
        RECT 159.800 95.200 160.100 128.800 ;
        RECT 160.600 126.800 161.000 127.200 ;
        RECT 163.000 126.800 163.400 127.200 ;
        RECT 160.600 125.200 160.900 126.800 ;
        RECT 163.000 126.200 163.300 126.800 ;
        RECT 161.400 126.100 161.800 126.200 ;
        RECT 162.200 126.100 162.600 126.200 ;
        RECT 161.400 125.800 162.600 126.100 ;
        RECT 163.000 125.800 163.400 126.200 ;
        RECT 163.800 125.200 164.100 135.800 ;
        RECT 164.600 135.100 165.000 135.200 ;
        RECT 165.400 135.100 165.800 135.200 ;
        RECT 164.600 134.800 165.800 135.100 ;
        RECT 166.200 134.800 166.600 135.200 ;
        RECT 168.600 135.100 169.000 135.200 ;
        RECT 169.400 135.100 169.800 135.200 ;
        RECT 168.600 134.800 169.800 135.100 ;
        RECT 166.200 134.200 166.500 134.800 ;
        RECT 164.600 133.800 165.000 134.200 ;
        RECT 165.400 134.100 165.800 134.200 ;
        RECT 166.200 134.100 166.600 134.200 ;
        RECT 165.400 133.800 166.600 134.100 ;
        RECT 167.000 134.100 167.400 134.200 ;
        RECT 167.800 134.100 168.200 134.200 ;
        RECT 167.000 133.800 168.200 134.100 ;
        RECT 168.600 133.800 169.000 134.200 ;
        RECT 164.600 133.200 164.900 133.800 ;
        RECT 164.600 132.800 165.000 133.200 ;
        RECT 166.200 127.200 166.500 133.800 ;
        RECT 167.000 132.800 167.400 133.200 ;
        RECT 167.000 132.200 167.300 132.800 ;
        RECT 167.000 131.800 167.400 132.200 ;
        RECT 168.600 129.200 168.900 133.800 ;
        RECT 170.200 133.100 170.600 135.900 ;
        RECT 171.800 132.100 172.200 137.900 ;
        RECT 175.800 135.200 176.100 146.800 ;
        RECT 179.000 143.100 179.400 148.900 ;
        RECT 182.200 148.800 182.600 149.200 ;
        RECT 182.200 145.100 182.600 147.900 ;
        RECT 183.000 147.200 183.300 151.800 ;
        RECT 183.000 146.800 183.400 147.200 ;
        RECT 180.600 143.100 181.000 143.200 ;
        RECT 181.400 143.100 181.800 143.200 ;
        RECT 180.600 142.800 181.800 143.100 ;
        RECT 172.600 134.700 173.000 135.200 ;
        RECT 175.800 134.800 176.200 135.200 ;
        RECT 172.600 134.200 172.900 134.700 ;
        RECT 172.600 133.800 173.000 134.200 ;
        RECT 168.600 128.800 169.000 129.200 ;
        RECT 167.000 127.800 167.400 128.200 ;
        RECT 167.000 127.200 167.300 127.800 ;
        RECT 167.800 127.500 168.200 127.900 ;
        RECT 168.500 127.500 170.600 127.800 ;
        RECT 171.100 127.500 171.500 127.900 ;
        RECT 166.200 126.800 166.600 127.200 ;
        RECT 167.000 126.800 167.400 127.200 ;
        RECT 167.800 127.100 168.100 127.500 ;
        RECT 168.500 127.400 168.900 127.500 ;
        RECT 170.200 127.400 170.600 127.500 ;
        RECT 167.800 126.800 170.200 127.100 ;
        RECT 165.400 125.800 165.800 126.200 ;
        RECT 160.600 124.800 161.000 125.200 ;
        RECT 163.800 124.800 164.200 125.200 ;
        RECT 160.600 108.200 160.900 124.800 ;
        RECT 163.800 119.200 164.100 124.800 ;
        RECT 165.400 122.200 165.700 125.800 ;
        RECT 167.800 125.100 168.100 126.800 ;
        RECT 169.800 126.700 170.200 126.800 ;
        RECT 171.200 125.100 171.500 127.500 ;
        RECT 167.800 124.700 168.200 125.100 ;
        RECT 171.100 124.700 171.500 125.100 ;
        RECT 171.800 126.800 172.200 127.200 ;
        RECT 171.800 125.200 172.100 126.800 ;
        RECT 171.800 124.800 172.200 125.200 ;
        RECT 171.800 123.800 172.200 124.200 ;
        RECT 174.200 123.800 174.600 124.200 ;
        RECT 165.400 121.800 165.800 122.200 ;
        RECT 163.800 118.800 164.200 119.200 ;
        RECT 161.400 112.100 161.800 117.900 ;
        RECT 164.600 115.000 165.000 115.100 ;
        RECT 165.400 115.000 165.800 115.100 ;
        RECT 164.600 114.700 165.800 115.000 ;
        RECT 164.600 112.200 164.900 114.700 ;
        RECT 164.600 111.800 165.000 112.200 ;
        RECT 166.200 112.100 166.600 117.900 ;
        RECT 168.600 116.800 169.000 117.200 ;
        RECT 168.600 116.200 168.900 116.800 ;
        RECT 167.000 113.800 167.400 114.200 ;
        RECT 167.000 113.200 167.300 113.800 ;
        RECT 167.000 112.800 167.400 113.200 ;
        RECT 167.800 113.100 168.200 115.900 ;
        RECT 168.600 115.800 169.000 116.200 ;
        RECT 169.400 112.800 169.800 113.200 ;
        RECT 162.200 109.800 162.600 110.200 ;
        RECT 162.200 108.200 162.500 109.800 ;
        RECT 164.600 108.800 165.000 109.200 ;
        RECT 160.600 107.800 161.000 108.200 ;
        RECT 162.200 108.100 162.600 108.200 ;
        RECT 163.000 108.100 163.400 108.200 ;
        RECT 162.200 107.800 163.400 108.100 ;
        RECT 160.600 106.200 160.900 107.800 ;
        RECT 164.600 107.200 164.900 108.800 ;
        RECT 167.000 107.800 167.400 108.200 ;
        RECT 167.000 107.200 167.300 107.800 ;
        RECT 161.400 107.100 161.800 107.200 ;
        RECT 162.200 107.100 162.600 107.200 ;
        RECT 161.400 106.800 162.600 107.100 ;
        RECT 164.600 106.800 165.000 107.200 ;
        RECT 167.000 107.100 167.400 107.200 ;
        RECT 167.800 107.100 168.200 107.200 ;
        RECT 167.000 106.800 168.200 107.100 ;
        RECT 168.600 106.800 169.000 107.200 ;
        RECT 168.600 106.200 168.900 106.800 ;
        RECT 160.600 105.800 161.000 106.200 ;
        RECT 163.000 106.100 163.400 106.200 ;
        RECT 163.800 106.100 164.200 106.200 ;
        RECT 163.000 105.800 164.200 106.100 ;
        RECT 165.400 106.100 165.800 106.200 ;
        RECT 166.200 106.100 166.600 106.200 ;
        RECT 165.400 105.800 166.600 106.100 ;
        RECT 167.800 105.800 168.200 106.200 ;
        RECT 168.600 105.800 169.000 106.200 ;
        RECT 159.800 94.800 160.200 95.200 ;
        RECT 161.400 92.100 161.800 97.900 ;
        RECT 163.000 93.100 163.400 95.900 ;
        RECT 163.800 93.100 164.200 95.900 ;
        RECT 165.400 92.100 165.800 97.900 ;
        RECT 166.200 94.700 166.600 95.100 ;
        RECT 166.200 94.200 166.500 94.700 ;
        RECT 166.200 93.800 166.600 94.200 ;
        RECT 167.800 91.200 168.100 105.800 ;
        RECT 169.400 95.200 169.700 112.800 ;
        RECT 171.000 112.100 171.400 117.900 ;
        RECT 171.800 111.200 172.100 123.800 ;
        RECT 172.600 121.800 173.000 122.200 ;
        RECT 172.600 116.200 172.900 121.800 ;
        RECT 172.600 115.800 173.000 116.200 ;
        RECT 173.400 114.800 173.800 115.200 ;
        RECT 171.800 110.800 172.200 111.200 ;
        RECT 171.800 106.200 172.100 110.800 ;
        RECT 173.400 109.200 173.700 114.800 ;
        RECT 174.200 114.200 174.500 123.800 ;
        RECT 175.000 123.100 175.400 128.900 ;
        RECT 175.800 126.200 176.100 134.800 ;
        RECT 176.600 132.100 177.000 137.900 ;
        RECT 180.600 133.800 181.000 134.200 ;
        RECT 179.000 131.800 179.400 132.200 ;
        RECT 175.800 125.800 176.200 126.200 ;
        RECT 177.400 126.100 177.800 126.200 ;
        RECT 178.200 126.100 178.600 126.200 ;
        RECT 177.400 125.800 178.600 126.100 ;
        RECT 175.000 116.800 175.400 117.200 ;
        RECT 175.000 115.100 175.300 116.800 ;
        RECT 175.000 114.700 175.400 115.100 ;
        RECT 174.200 113.800 174.600 114.200 ;
        RECT 173.400 108.800 173.800 109.200 ;
        RECT 174.200 108.200 174.500 113.800 ;
        RECT 175.800 112.100 176.200 117.900 ;
        RECT 177.400 117.200 177.700 125.800 ;
        RECT 179.000 125.200 179.300 131.800 ;
        RECT 179.000 124.800 179.400 125.200 ;
        RECT 179.800 123.100 180.200 128.900 ;
        RECT 179.000 121.800 179.400 122.200 ;
        RECT 177.400 116.800 177.800 117.200 ;
        RECT 176.600 113.800 177.000 114.200 ;
        RECT 176.600 113.200 176.900 113.800 ;
        RECT 176.600 112.800 177.000 113.200 ;
        RECT 177.400 113.100 177.800 115.900 ;
        RECT 179.000 115.200 179.300 121.800 ;
        RECT 179.800 115.800 180.200 116.200 ;
        RECT 179.800 115.200 180.100 115.800 ;
        RECT 179.000 114.800 179.400 115.200 ;
        RECT 179.800 114.800 180.200 115.200 ;
        RECT 180.600 113.200 180.900 133.800 ;
        RECT 182.200 132.100 182.600 137.900 ;
        RECT 183.000 135.200 183.300 146.800 ;
        RECT 183.800 143.100 184.200 148.900 ;
        RECT 184.600 145.900 185.000 146.300 ;
        RECT 184.600 145.200 184.900 145.900 ;
        RECT 184.600 144.800 185.000 145.200 ;
        RECT 188.600 143.100 189.000 148.900 ;
        RECT 190.200 143.100 190.600 143.200 ;
        RECT 191.000 143.100 191.400 143.200 ;
        RECT 190.200 142.800 191.400 143.100 ;
        RECT 183.000 134.800 183.400 135.200 ;
        RECT 183.800 135.100 184.200 135.200 ;
        RECT 184.600 135.100 185.000 135.200 ;
        RECT 183.800 134.800 185.000 135.100 ;
        RECT 183.000 134.200 183.300 134.800 ;
        RECT 183.000 133.800 183.400 134.200 ;
        RECT 187.000 132.100 187.400 137.900 ;
        RECT 188.600 133.100 189.000 135.900 ;
        RECT 191.800 134.800 192.200 135.200 ;
        RECT 188.600 128.800 189.000 129.200 ;
        RECT 188.600 128.200 188.900 128.800 ;
        RECT 183.800 128.100 184.200 128.200 ;
        RECT 184.600 128.100 185.000 128.200 ;
        RECT 181.400 125.100 181.800 127.900 ;
        RECT 183.800 127.800 185.000 128.100 ;
        RECT 187.000 127.800 187.400 128.200 ;
        RECT 188.600 127.800 189.000 128.200 ;
        RECT 183.000 125.800 183.400 126.200 ;
        RECT 186.200 126.100 186.600 126.200 ;
        RECT 187.000 126.100 187.300 127.800 ;
        RECT 191.800 127.200 192.100 134.800 ;
        RECT 193.400 127.800 193.800 128.200 ;
        RECT 191.800 126.800 192.200 127.200 ;
        RECT 186.200 125.800 187.300 126.100 ;
        RECT 188.600 126.100 189.000 126.200 ;
        RECT 189.400 126.100 189.800 126.200 ;
        RECT 188.600 125.800 189.800 126.100 ;
        RECT 190.200 125.800 190.600 126.200 ;
        RECT 191.000 126.100 191.400 126.200 ;
        RECT 191.800 126.100 192.200 126.200 ;
        RECT 191.000 125.800 192.200 126.100 ;
        RECT 183.000 124.200 183.300 125.800 ;
        RECT 183.000 123.800 183.400 124.200 ;
        RECT 186.200 118.200 186.500 125.800 ;
        RECT 189.400 123.800 189.800 124.200 ;
        RECT 182.200 117.800 182.600 118.200 ;
        RECT 186.200 118.100 186.600 118.200 ;
        RECT 186.200 117.800 187.300 118.100 ;
        RECT 182.200 115.200 182.500 117.800 ;
        RECT 183.000 115.800 183.400 116.200 ;
        RECT 183.800 115.800 184.200 116.200 ;
        RECT 186.200 115.800 186.600 116.200 ;
        RECT 183.000 115.200 183.300 115.800 ;
        RECT 183.800 115.200 184.100 115.800 ;
        RECT 186.200 115.200 186.500 115.800 ;
        RECT 182.200 114.800 182.600 115.200 ;
        RECT 183.000 114.800 183.400 115.200 ;
        RECT 183.800 114.800 184.200 115.200 ;
        RECT 184.600 115.100 185.000 115.200 ;
        RECT 185.400 115.100 185.800 115.200 ;
        RECT 184.600 114.800 185.800 115.100 ;
        RECT 186.200 114.800 186.600 115.200 ;
        RECT 185.400 114.100 185.800 114.200 ;
        RECT 184.600 113.800 185.800 114.100 ;
        RECT 180.600 112.800 181.000 113.200 ;
        RECT 180.600 109.200 180.900 112.800 ;
        RECT 184.600 109.200 184.900 113.800 ;
        RECT 185.400 113.200 185.700 113.800 ;
        RECT 185.400 112.800 185.800 113.200 ;
        RECT 180.600 108.800 181.000 109.200 ;
        RECT 184.600 108.800 185.000 109.200 ;
        RECT 174.200 107.800 174.600 108.200 ;
        RECT 171.800 105.800 172.200 106.200 ;
        RECT 169.400 94.800 169.800 95.200 ;
        RECT 169.400 93.800 169.800 94.200 ;
        RECT 167.800 90.800 168.200 91.200 ;
        RECT 159.800 89.800 160.200 90.200 ;
        RECT 159.800 89.200 160.100 89.800 ;
        RECT 150.200 86.800 150.600 87.200 ;
        RECT 151.000 86.800 151.400 87.200 ;
        RECT 150.200 86.200 150.500 86.800 ;
        RECT 150.200 85.800 150.600 86.200 ;
        RECT 152.600 83.100 153.000 88.900 ;
        RECT 159.800 88.800 160.200 89.200 ;
        RECT 169.400 88.200 169.700 93.800 ;
        RECT 170.200 92.100 170.600 97.900 ;
        RECT 172.600 96.800 173.000 97.200 ;
        RECT 172.600 94.200 172.900 96.800 ;
        RECT 174.200 95.200 174.500 107.800 ;
        RECT 187.000 106.200 187.300 117.800 ;
        RECT 189.400 115.200 189.700 123.800 ;
        RECT 190.200 115.200 190.500 125.800 ;
        RECT 193.400 124.200 193.700 127.800 ;
        RECT 193.400 123.800 193.800 124.200 ;
        RECT 188.600 114.800 189.000 115.200 ;
        RECT 189.400 114.800 189.800 115.200 ;
        RECT 190.200 114.800 190.600 115.200 ;
        RECT 188.600 114.200 188.900 114.800 ;
        RECT 189.400 114.200 189.700 114.800 ;
        RECT 188.600 113.800 189.000 114.200 ;
        RECT 189.400 113.800 189.800 114.200 ;
        RECT 189.400 109.200 189.700 113.800 ;
        RECT 190.200 113.100 190.600 113.200 ;
        RECT 191.000 113.100 191.400 113.200 ;
        RECT 190.200 112.800 191.400 113.100 ;
        RECT 194.200 109.200 194.500 161.800 ;
        RECT 195.000 126.800 195.400 127.200 ;
        RECT 195.000 126.200 195.300 126.800 ;
        RECT 195.000 125.800 195.400 126.200 ;
        RECT 195.000 121.800 195.400 122.200 ;
        RECT 189.400 108.800 189.800 109.200 ;
        RECT 191.800 108.800 192.200 109.200 ;
        RECT 194.200 108.800 194.600 109.200 ;
        RECT 191.800 108.200 192.100 108.800 ;
        RECT 191.800 107.800 192.200 108.200 ;
        RECT 190.200 106.800 190.600 107.200 ;
        RECT 190.200 106.200 190.500 106.800 ;
        RECT 182.200 106.100 182.600 106.200 ;
        RECT 183.000 106.100 183.400 106.200 ;
        RECT 182.200 105.800 183.400 106.100 ;
        RECT 187.000 105.800 187.400 106.200 ;
        RECT 190.200 105.800 190.600 106.200 ;
        RECT 180.600 101.800 181.000 102.200 ;
        RECT 180.600 99.200 180.900 101.800 ;
        RECT 180.600 98.800 181.000 99.200 ;
        RECT 183.800 98.800 184.200 99.200 ;
        RECT 174.200 94.800 174.600 95.200 ;
        RECT 172.600 93.800 173.000 94.200 ;
        RECT 171.800 91.800 172.200 92.200 ;
        RECT 172.600 92.100 173.000 92.200 ;
        RECT 173.400 92.100 173.800 92.200 ;
        RECT 175.800 92.100 176.200 97.900 ;
        RECT 176.600 95.800 177.000 96.200 ;
        RECT 176.600 95.200 176.900 95.800 ;
        RECT 176.600 94.800 177.000 95.200 ;
        RECT 179.000 94.800 179.400 95.200 ;
        RECT 172.600 91.800 173.800 92.100 ;
        RECT 153.400 86.800 153.800 87.200 ;
        RECT 153.400 79.200 153.700 86.800 ;
        RECT 154.200 85.100 154.600 87.900 ;
        RECT 169.400 87.800 169.800 88.200 ;
        RECT 169.400 87.200 169.700 87.800 ;
        RECT 171.800 87.200 172.100 91.800 ;
        RECT 179.000 88.200 179.300 94.800 ;
        RECT 180.600 92.100 181.000 97.900 ;
        RECT 182.200 93.100 182.600 95.900 ;
        RECT 183.000 93.100 183.400 95.900 ;
        RECT 183.800 94.200 184.100 98.800 ;
        RECT 183.800 93.800 184.200 94.200 ;
        RECT 183.800 89.200 184.100 93.800 ;
        RECT 184.600 92.100 185.000 97.900 ;
        RECT 185.400 95.000 185.800 95.100 ;
        RECT 186.200 95.000 186.600 95.100 ;
        RECT 185.400 94.700 186.600 95.000 ;
        RECT 189.400 92.100 189.800 97.900 ;
        RECT 191.000 92.100 191.400 92.200 ;
        RECT 191.800 92.100 192.200 92.200 ;
        RECT 191.000 91.800 192.200 92.100 ;
        RECT 195.000 91.200 195.300 121.800 ;
        RECT 191.800 90.800 192.200 91.200 ;
        RECT 195.000 90.800 195.400 91.200 ;
        RECT 183.800 88.800 184.200 89.200 ;
        RECT 174.200 87.800 174.600 88.200 ;
        RECT 175.800 88.100 176.200 88.200 ;
        RECT 176.600 88.100 177.000 88.200 ;
        RECT 175.800 87.800 177.000 88.100 ;
        RECT 179.000 87.800 179.400 88.200 ;
        RECT 181.400 87.800 181.800 88.200 ;
        RECT 157.400 86.800 157.800 87.200 ;
        RECT 162.200 86.800 162.600 87.200 ;
        RECT 163.800 87.100 164.200 87.200 ;
        RECT 163.000 86.800 164.200 87.100 ;
        RECT 169.400 86.800 169.800 87.200 ;
        RECT 171.800 86.800 172.200 87.200 ;
        RECT 173.400 86.800 173.800 87.200 ;
        RECT 157.400 86.200 157.700 86.800 ;
        RECT 157.400 85.800 157.800 86.200 ;
        RECT 162.200 82.200 162.500 86.800 ;
        RECT 162.200 81.800 162.600 82.200 ;
        RECT 163.000 79.200 163.300 86.800 ;
        RECT 163.800 84.200 164.100 86.800 ;
        RECT 164.600 86.100 165.000 86.200 ;
        RECT 165.400 86.100 165.800 86.200 ;
        RECT 164.600 85.800 165.800 86.100 ;
        RECT 166.200 85.800 166.600 86.200 ;
        RECT 167.800 85.800 168.200 86.200 ;
        RECT 166.200 85.200 166.500 85.800 ;
        RECT 167.800 85.200 168.100 85.800 ;
        RECT 165.400 84.800 165.800 85.200 ;
        RECT 166.200 84.800 166.600 85.200 ;
        RECT 167.800 84.800 168.200 85.200 ;
        RECT 163.800 83.800 164.200 84.200 ;
        RECT 164.600 82.800 165.000 83.200 ;
        RECT 164.600 82.200 164.900 82.800 ;
        RECT 165.400 82.200 165.700 84.800 ;
        RECT 164.600 81.800 165.000 82.200 ;
        RECT 165.400 81.800 165.800 82.200 ;
        RECT 137.400 78.800 137.800 79.200 ;
        RECT 153.400 78.800 153.800 79.200 ;
        RECT 163.000 78.800 163.400 79.200 ;
        RECT 137.400 78.200 137.700 78.800 ;
        RECT 137.400 77.800 137.800 78.200 ;
        RECT 134.200 74.100 134.600 74.200 ;
        RECT 135.000 74.100 135.400 74.200 ;
        RECT 134.200 73.800 135.400 74.100 ;
        RECT 136.600 73.800 137.000 74.200 ;
        RECT 137.400 74.100 137.800 74.200 ;
        RECT 138.200 74.100 138.600 74.200 ;
        RECT 137.400 73.800 138.600 74.100 ;
        RECT 139.000 73.100 139.400 75.900 ;
        RECT 140.600 72.100 141.000 77.900 ;
        RECT 142.200 74.800 142.600 75.200 ;
        RECT 139.800 69.800 140.200 70.200 ;
        RECT 139.800 69.200 140.100 69.800 ;
        RECT 131.000 65.100 131.400 67.900 ;
        RECT 122.200 64.100 122.600 64.200 ;
        RECT 123.000 64.100 123.400 64.200 ;
        RECT 122.200 63.800 123.400 64.100 ;
        RECT 124.600 63.800 125.000 64.200 ;
        RECT 132.600 63.100 133.000 68.900 ;
        RECT 133.400 68.800 133.800 69.200 ;
        RECT 133.400 68.200 133.700 68.800 ;
        RECT 133.400 67.800 133.800 68.200 ;
        RECT 134.200 66.100 134.600 66.200 ;
        RECT 135.000 66.100 135.400 66.200 ;
        RECT 134.200 65.800 135.400 66.100 ;
        RECT 137.400 63.100 137.800 68.900 ;
        RECT 139.800 68.800 140.200 69.200 ;
        RECT 142.200 66.200 142.500 74.800 ;
        RECT 145.400 72.100 145.800 77.900 ;
        RECT 146.200 73.800 146.600 74.200 ;
        RECT 146.200 69.200 146.500 73.800 ;
        RECT 152.600 72.800 153.000 73.200 ;
        RECT 154.200 73.100 154.600 75.900 ;
        RECT 155.000 73.800 155.400 74.200 ;
        RECT 155.000 73.200 155.300 73.800 ;
        RECT 155.000 72.800 155.400 73.200 ;
        RECT 152.600 72.200 152.900 72.800 ;
        RECT 147.800 71.800 148.200 72.200 ;
        RECT 152.600 71.800 153.000 72.200 ;
        RECT 147.800 70.200 148.100 71.800 ;
        RECT 147.800 69.800 148.200 70.200 ;
        RECT 155.000 69.200 155.300 72.800 ;
        RECT 155.800 72.100 156.200 77.900 ;
        RECT 158.200 75.100 158.600 75.200 ;
        RECT 159.000 75.100 159.400 75.200 ;
        RECT 158.200 74.800 159.400 75.100 ;
        RECT 160.600 72.100 161.000 77.900 ;
        RECT 164.600 76.200 164.900 81.800 ;
        RECT 166.200 77.200 166.500 84.800 ;
        RECT 167.800 84.100 168.200 84.200 ;
        RECT 168.600 84.100 169.000 84.200 ;
        RECT 167.800 83.800 169.000 84.100 ;
        RECT 170.200 84.100 170.600 84.200 ;
        RECT 171.000 84.100 171.400 84.200 ;
        RECT 170.200 83.800 171.400 84.100 ;
        RECT 173.400 83.200 173.700 86.800 ;
        RECT 174.200 86.200 174.500 87.800 ;
        RECT 181.400 87.200 181.700 87.800 ;
        RECT 182.200 87.500 182.600 87.900 ;
        RECT 182.900 87.500 185.000 87.800 ;
        RECT 185.500 87.500 185.900 87.900 ;
        RECT 181.400 86.800 181.800 87.200 ;
        RECT 182.200 87.100 182.500 87.500 ;
        RECT 182.900 87.400 183.300 87.500 ;
        RECT 184.600 87.400 185.000 87.500 ;
        RECT 182.200 86.800 184.600 87.100 ;
        RECT 174.200 85.800 174.600 86.200 ;
        RECT 178.200 85.800 178.600 86.200 ;
        RECT 179.000 85.800 179.400 86.200 ;
        RECT 175.000 85.100 175.400 85.200 ;
        RECT 175.800 85.100 176.200 85.200 ;
        RECT 175.000 84.800 176.200 85.100 ;
        RECT 178.200 83.200 178.500 85.800 ;
        RECT 173.400 82.800 173.800 83.200 ;
        RECT 178.200 82.800 178.600 83.200 ;
        RECT 167.000 81.800 167.400 82.200 ;
        RECT 174.200 81.800 174.600 82.200 ;
        RECT 178.200 81.800 178.600 82.200 ;
        RECT 166.200 76.800 166.600 77.200 ;
        RECT 164.600 75.800 165.000 76.200 ;
        RECT 166.200 75.800 166.600 76.200 ;
        RECT 163.800 74.800 164.200 75.200 ;
        RECT 164.600 75.100 165.000 75.200 ;
        RECT 165.400 75.100 165.800 75.200 ;
        RECT 164.600 74.800 165.800 75.100 ;
        RECT 163.000 73.800 163.400 74.200 ;
        RECT 163.000 73.200 163.300 73.800 ;
        RECT 163.000 72.800 163.400 73.200 ;
        RECT 163.800 71.200 164.100 74.800 ;
        RECT 166.200 74.200 166.500 75.800 ;
        RECT 167.000 74.200 167.300 81.800 ;
        RECT 173.400 76.800 173.800 77.200 ;
        RECT 167.800 76.100 168.200 76.200 ;
        RECT 168.600 76.100 169.000 76.200 ;
        RECT 167.800 75.800 169.000 76.100 ;
        RECT 170.200 75.800 170.600 76.200 ;
        RECT 170.200 75.200 170.500 75.800 ;
        RECT 170.200 74.800 170.600 75.200 ;
        RECT 164.600 73.800 165.000 74.200 ;
        RECT 166.200 73.800 166.600 74.200 ;
        RECT 167.000 73.800 167.400 74.200 ;
        RECT 172.600 74.100 173.000 74.200 ;
        RECT 171.800 73.800 173.000 74.100 ;
        RECT 163.800 70.800 164.200 71.200 ;
        RECT 163.800 69.200 164.100 70.800 ;
        RECT 146.200 68.800 146.600 69.200 ;
        RECT 155.000 68.800 155.400 69.200 ;
        RECT 163.800 68.800 164.200 69.200 ;
        RECT 160.600 67.800 161.000 68.200 ;
        RECT 160.600 67.200 160.900 67.800 ;
        RECT 164.600 67.200 164.900 73.800 ;
        RECT 165.400 72.800 165.800 73.200 ;
        RECT 168.600 73.100 169.000 73.200 ;
        RECT 169.400 73.100 169.800 73.200 ;
        RECT 168.600 72.800 169.800 73.100 ;
        RECT 165.400 72.200 165.700 72.800 ;
        RECT 165.400 71.800 165.800 72.200 ;
        RECT 167.000 72.100 167.400 72.200 ;
        RECT 167.800 72.100 168.200 72.200 ;
        RECT 167.000 71.800 168.200 72.100 ;
        RECT 166.200 68.800 166.600 69.200 ;
        RECT 166.200 67.200 166.500 68.800 ;
        RECT 171.800 68.200 172.100 73.800 ;
        RECT 169.400 67.800 169.800 68.200 ;
        RECT 171.800 67.800 172.200 68.200 ;
        RECT 169.400 67.200 169.700 67.800 ;
        RECT 154.200 67.100 154.600 67.200 ;
        RECT 155.000 67.100 155.400 67.200 ;
        RECT 154.200 66.800 155.400 67.100 ;
        RECT 159.000 66.800 159.400 67.200 ;
        RECT 159.800 66.800 160.200 67.200 ;
        RECT 160.600 66.800 161.000 67.200 ;
        RECT 162.200 67.100 162.600 67.200 ;
        RECT 163.000 67.100 163.400 67.200 ;
        RECT 162.200 66.800 163.400 67.100 ;
        RECT 164.600 66.800 165.000 67.200 ;
        RECT 166.200 66.800 166.600 67.200 ;
        RECT 169.400 66.800 169.800 67.200 ;
        RECT 170.200 66.800 170.600 67.200 ;
        RECT 159.000 66.200 159.300 66.800 ;
        RECT 142.200 65.800 142.600 66.200 ;
        RECT 147.000 65.800 147.400 66.200 ;
        RECT 153.400 66.100 153.800 66.200 ;
        RECT 154.200 66.100 154.600 66.200 ;
        RECT 155.000 66.100 155.400 66.200 ;
        RECT 153.400 65.800 155.400 66.100 ;
        RECT 159.000 65.800 159.400 66.200 ;
        RECT 129.400 61.800 129.800 62.200 ;
        RECT 139.800 61.800 140.200 62.200 ;
        RECT 111.000 58.800 111.400 59.200 ;
        RECT 105.400 56.800 105.800 57.200 ;
        RECT 110.200 56.800 110.600 57.200 ;
        RECT 115.800 56.800 116.200 57.200 ;
        RECT 80.600 55.800 81.000 56.200 ;
        RECT 83.000 56.100 83.400 56.200 ;
        RECT 83.800 56.100 84.200 56.200 ;
        RECT 83.000 55.800 84.200 56.100 ;
        RECT 86.200 55.800 86.600 56.200 ;
        RECT 87.000 55.800 87.400 56.200 ;
        RECT 103.800 55.800 104.200 56.200 ;
        RECT 105.400 55.800 105.800 56.200 ;
        RECT 80.600 55.200 80.900 55.800 ;
        RECT 71.000 54.800 71.400 55.200 ;
        RECT 72.600 54.800 73.000 55.200 ;
        RECT 75.000 54.800 75.400 55.200 ;
        RECT 75.800 54.800 76.200 55.200 ;
        RECT 76.600 54.800 77.000 55.200 ;
        RECT 79.000 54.800 79.400 55.200 ;
        RECT 80.600 54.800 81.000 55.200 ;
        RECT 83.800 54.800 84.200 55.200 ;
        RECT 71.000 54.200 71.300 54.800 ;
        RECT 72.600 54.200 72.900 54.800 ;
        RECT 83.800 54.200 84.100 54.800 ;
        RECT 86.200 54.200 86.500 55.800 ;
        RECT 87.000 55.200 87.300 55.800 ;
        RECT 103.800 55.200 104.100 55.800 ;
        RECT 105.400 55.200 105.700 55.800 ;
        RECT 87.000 54.800 87.400 55.200 ;
        RECT 87.800 55.100 88.200 55.200 ;
        RECT 88.600 55.100 89.000 55.200 ;
        RECT 87.800 54.800 89.000 55.100 ;
        RECT 103.800 54.800 104.200 55.200 ;
        RECT 105.400 54.800 105.800 55.200 ;
        RECT 106.200 54.800 106.600 55.200 ;
        RECT 107.800 55.100 108.200 55.200 ;
        RECT 108.600 55.100 109.000 55.200 ;
        RECT 107.800 54.800 109.000 55.100 ;
        RECT 109.400 54.800 109.800 55.200 ;
        RECT 71.000 53.800 71.400 54.200 ;
        RECT 72.600 53.800 73.000 54.200 ;
        RECT 77.400 53.800 77.800 54.200 ;
        RECT 83.800 53.800 84.200 54.200 ;
        RECT 86.200 53.800 86.600 54.200 ;
        RECT 87.800 53.800 88.200 54.200 ;
        RECT 90.200 53.800 90.600 54.200 ;
        RECT 95.800 53.800 96.200 54.200 ;
        RECT 103.000 53.800 103.400 54.200 ;
        RECT 77.400 53.200 77.700 53.800 ;
        RECT 87.800 53.200 88.100 53.800 ;
        RECT 90.200 53.200 90.500 53.800 ;
        RECT 71.000 52.800 71.400 53.200 ;
        RECT 72.600 53.100 73.000 53.200 ;
        RECT 73.400 53.100 73.800 53.200 ;
        RECT 72.600 52.800 73.800 53.100 ;
        RECT 77.400 52.800 77.800 53.200 ;
        RECT 83.800 53.100 84.200 53.200 ;
        RECT 84.600 53.100 85.000 53.200 ;
        RECT 83.800 52.800 85.000 53.100 ;
        RECT 86.200 52.800 86.600 53.200 ;
        RECT 87.000 53.100 87.400 53.200 ;
        RECT 87.800 53.100 88.200 53.200 ;
        RECT 87.000 52.800 88.200 53.100 ;
        RECT 90.200 52.800 90.600 53.200 ;
        RECT 92.600 53.100 93.000 53.200 ;
        RECT 91.800 52.800 93.000 53.100 ;
        RECT 93.400 52.800 93.800 53.200 ;
        RECT 95.000 52.800 95.400 53.200 ;
        RECT 71.000 52.200 71.300 52.800 ;
        RECT 71.000 51.800 71.400 52.200 ;
        RECT 68.600 48.800 69.700 49.100 ;
        RECT 67.800 48.100 68.200 48.200 ;
        RECT 68.600 48.100 69.000 48.200 ;
        RECT 67.800 47.800 69.000 48.100 ;
        RECT 71.000 43.100 71.400 48.900 ;
        RECT 73.400 47.200 73.700 52.800 ;
        RECT 74.200 51.800 74.600 52.200 ;
        RECT 73.400 46.800 73.800 47.200 ;
        RECT 74.200 46.200 74.500 51.800 ;
        RECT 78.200 49.100 78.600 49.200 ;
        RECT 79.000 49.100 79.400 49.200 ;
        RECT 74.200 45.800 74.600 46.200 ;
        RECT 75.800 43.100 76.200 48.900 ;
        RECT 78.200 48.800 79.400 49.100 ;
        RECT 77.400 45.100 77.800 47.900 ;
        RECT 80.600 47.800 81.000 48.200 ;
        RECT 83.000 47.800 83.400 48.200 ;
        RECT 80.600 47.200 80.900 47.800 ;
        RECT 80.600 46.800 81.000 47.200 ;
        RECT 81.400 47.100 81.800 47.200 ;
        RECT 82.200 47.100 82.600 47.200 ;
        RECT 81.400 46.800 82.600 47.100 ;
        RECT 83.000 45.200 83.300 47.800 ;
        RECT 78.200 44.800 78.600 45.200 ;
        RECT 83.000 44.800 83.400 45.200 ;
        RECT 59.800 34.700 60.200 35.100 ;
        RECT 47.800 29.100 48.200 29.200 ;
        RECT 48.600 29.100 49.000 29.200 ;
        RECT 42.200 25.900 42.600 26.300 ;
        RECT 46.200 23.100 46.600 28.900 ;
        RECT 47.800 28.800 49.000 29.100 ;
        RECT 54.200 28.800 54.600 29.200 ;
        RECT 51.000 26.800 51.400 27.200 ;
        RECT 51.000 24.200 51.300 26.800 ;
        RECT 51.000 23.800 51.400 24.200 ;
        RECT 56.600 23.100 57.000 28.900 ;
        RECT 59.800 28.100 60.100 34.700 ;
        RECT 60.600 32.100 61.000 37.900 ;
        RECT 78.200 37.200 78.500 44.800 ;
        RECT 78.200 36.800 78.600 37.200 ;
        RECT 61.400 33.800 61.800 34.200 ;
        RECT 61.400 32.100 61.700 33.800 ;
        RECT 62.200 33.100 62.600 35.900 ;
        RECT 69.400 35.800 69.800 36.200 ;
        RECT 69.400 35.200 69.700 35.800 ;
        RECT 67.800 34.800 68.200 35.200 ;
        RECT 69.400 34.800 69.800 35.200 ;
        RECT 67.800 34.200 68.100 34.800 ;
        RECT 67.800 33.800 68.200 34.200 ;
        RECT 71.800 34.100 72.200 34.200 ;
        RECT 72.600 34.100 73.000 34.200 ;
        RECT 71.800 33.800 73.000 34.100 ;
        RECT 75.000 33.800 75.400 34.200 ;
        RECT 66.200 32.800 66.600 33.200 ;
        RECT 61.400 31.800 62.500 32.100 ;
        RECT 59.800 27.800 60.900 28.100 ;
        RECT 59.800 26.800 60.200 27.200 ;
        RECT 23.800 16.800 24.200 17.200 ;
        RECT 35.000 16.800 35.400 17.200 ;
        RECT 36.600 16.800 37.000 17.200 ;
        RECT 31.800 15.800 32.200 16.200 ;
        RECT 31.800 15.200 32.100 15.800 ;
        RECT 35.000 15.200 35.300 16.800 ;
        RECT 23.800 15.100 24.200 15.200 ;
        RECT 24.600 15.100 25.000 15.200 ;
        RECT 23.800 14.800 25.000 15.100 ;
        RECT 27.000 14.800 27.400 15.200 ;
        RECT 29.400 14.800 29.800 15.200 ;
        RECT 31.800 14.800 32.200 15.200 ;
        RECT 34.200 15.100 34.600 15.200 ;
        RECT 33.400 14.800 34.600 15.100 ;
        RECT 35.000 14.800 35.400 15.200 ;
        RECT 26.200 13.800 26.600 14.200 ;
        RECT 26.200 13.200 26.500 13.800 ;
        RECT 26.200 12.800 26.600 13.200 ;
        RECT 27.000 12.200 27.300 14.800 ;
        RECT 27.800 13.800 28.200 14.200 ;
        RECT 28.600 13.800 29.000 14.200 ;
        RECT 23.000 12.100 23.400 12.200 ;
        RECT 23.800 12.100 24.200 12.200 ;
        RECT 23.000 11.800 24.200 12.100 ;
        RECT 27.000 11.800 27.400 12.200 ;
        RECT 27.800 11.100 28.100 13.800 ;
        RECT 28.600 13.200 28.900 13.800 ;
        RECT 29.400 13.200 29.700 14.800 ;
        RECT 30.200 13.800 30.600 14.200 ;
        RECT 28.600 12.800 29.000 13.200 ;
        RECT 29.400 12.800 29.800 13.200 ;
        RECT 30.200 12.200 30.500 13.800 ;
        RECT 31.000 12.800 31.400 13.200 ;
        RECT 30.200 11.800 30.600 12.200 ;
        RECT 27.000 10.800 28.100 11.100 ;
        RECT 30.200 10.800 30.600 11.200 ;
        RECT 27.000 10.200 27.300 10.800 ;
        RECT 27.000 9.800 27.400 10.200 ;
        RECT 19.000 8.800 19.400 9.200 ;
        RECT 21.400 8.800 21.800 9.200 ;
        RECT 20.600 7.800 21.000 8.200 ;
        RECT 8.600 6.800 9.000 7.200 ;
        RECT 11.000 7.100 11.400 7.200 ;
        RECT 11.800 7.100 12.200 7.200 ;
        RECT 11.000 6.800 12.200 7.100 ;
        RECT 15.800 6.800 16.200 7.200 ;
        RECT 17.400 7.100 17.800 7.200 ;
        RECT 18.200 7.100 18.600 7.200 ;
        RECT 17.400 6.800 18.600 7.100 ;
        RECT 20.600 6.200 20.900 7.800 ;
        RECT 21.400 7.200 21.700 8.800 ;
        RECT 27.000 8.200 27.300 9.800 ;
        RECT 30.200 9.200 30.500 10.800 ;
        RECT 31.000 9.200 31.300 12.800 ;
        RECT 33.400 9.200 33.700 14.800 ;
        RECT 34.200 12.800 34.600 13.200 ;
        RECT 30.200 8.800 30.600 9.200 ;
        RECT 31.000 8.800 31.400 9.200 ;
        RECT 33.400 8.800 33.800 9.200 ;
        RECT 23.800 7.800 24.200 8.200 ;
        RECT 27.000 7.800 27.400 8.200 ;
        RECT 29.400 8.100 29.800 8.200 ;
        RECT 30.200 8.100 30.600 8.200 ;
        RECT 29.400 7.800 30.600 8.100 ;
        RECT 23.800 7.200 24.100 7.800 ;
        RECT 31.000 7.200 31.300 8.800 ;
        RECT 32.600 7.800 33.000 8.200 ;
        RECT 21.400 6.800 21.800 7.200 ;
        RECT 22.200 7.100 22.600 7.200 ;
        RECT 23.000 7.100 23.400 7.200 ;
        RECT 22.200 6.800 23.400 7.100 ;
        RECT 23.800 6.800 24.200 7.200 ;
        RECT 31.000 6.800 31.400 7.200 ;
        RECT 3.000 6.100 3.400 6.200 ;
        RECT 3.800 6.100 4.200 6.200 ;
        RECT 3.000 5.800 4.200 6.100 ;
        RECT 14.200 5.800 14.600 6.200 ;
        RECT 15.000 6.100 15.400 6.200 ;
        RECT 15.800 6.100 16.200 6.200 ;
        RECT 15.000 5.800 16.200 6.100 ;
        RECT 16.600 5.800 17.000 6.200 ;
        RECT 20.600 5.800 21.000 6.200 ;
        RECT 25.400 5.800 25.800 6.200 ;
        RECT 29.400 5.800 29.800 6.200 ;
        RECT 14.200 5.200 14.500 5.800 ;
        RECT 16.600 5.200 16.900 5.800 ;
        RECT 4.600 5.100 5.000 5.200 ;
        RECT 5.400 5.100 5.800 5.200 ;
        RECT 4.600 4.800 5.800 5.100 ;
        RECT 14.200 4.800 14.600 5.200 ;
        RECT 15.800 5.100 16.200 5.200 ;
        RECT 16.600 5.100 17.000 5.200 ;
        RECT 15.800 4.800 17.000 5.100 ;
        RECT 19.000 5.100 19.400 5.200 ;
        RECT 19.800 5.100 20.200 5.200 ;
        RECT 19.000 4.800 20.200 5.100 ;
        RECT 25.400 4.200 25.700 5.800 ;
        RECT 29.400 4.200 29.700 5.800 ;
        RECT 32.600 5.200 32.900 7.800 ;
        RECT 34.200 7.200 34.500 12.800 ;
        RECT 37.400 12.100 37.800 17.900 ;
        RECT 40.600 15.200 40.900 22.800 ;
        RECT 59.800 19.200 60.100 26.800 ;
        RECT 60.600 26.300 60.900 27.800 ;
        RECT 60.600 25.900 61.000 26.300 ;
        RECT 61.400 23.100 61.800 28.900 ;
        RECT 59.800 18.800 60.200 19.200 ;
        RECT 41.400 15.800 41.800 16.200 ;
        RECT 40.600 14.800 41.000 15.200 ;
        RECT 41.400 10.200 41.700 15.800 ;
        RECT 42.200 12.100 42.600 17.900 ;
        RECT 47.000 16.800 47.400 17.200 ;
        RECT 48.600 17.100 49.000 17.200 ;
        RECT 49.400 17.100 49.800 17.200 ;
        RECT 48.600 16.800 49.800 17.100 ;
        RECT 43.000 13.800 43.400 14.200 ;
        RECT 43.000 13.200 43.300 13.800 ;
        RECT 43.000 12.800 43.400 13.200 ;
        RECT 43.800 13.100 44.200 15.900 ;
        RECT 47.000 15.200 47.300 16.800 ;
        RECT 47.000 14.800 47.400 15.200 ;
        RECT 46.200 13.800 46.600 14.200 ;
        RECT 46.200 11.200 46.500 13.800 ;
        RECT 45.400 10.800 45.800 11.200 ;
        RECT 46.200 10.800 46.600 11.200 ;
        RECT 41.400 9.800 41.800 10.200 ;
        RECT 35.000 9.100 35.400 9.200 ;
        RECT 35.800 9.100 36.200 9.200 ;
        RECT 35.000 8.800 36.200 9.100 ;
        RECT 34.200 6.800 34.600 7.200 ;
        RECT 32.600 4.800 33.000 5.200 ;
        RECT 25.400 3.800 25.800 4.200 ;
        RECT 29.400 3.800 29.800 4.200 ;
        RECT 37.400 3.100 37.800 8.900 ;
        RECT 41.400 8.200 41.700 9.800 ;
        RECT 41.400 7.800 41.800 8.200 ;
        RECT 41.400 5.900 41.800 6.300 ;
        RECT 41.400 5.200 41.700 5.900 ;
        RECT 41.400 4.800 41.800 5.200 ;
        RECT 42.200 3.100 42.600 8.900 ;
        RECT 43.800 5.100 44.200 7.900 ;
        RECT 45.400 6.200 45.700 10.800 ;
        RECT 47.000 9.200 47.300 14.800 ;
        RECT 48.600 11.800 49.000 12.200 ;
        RECT 50.200 11.800 50.600 12.200 ;
        RECT 51.800 12.100 52.200 17.900 ;
        RECT 55.000 14.800 55.400 15.200 ;
        RECT 55.800 14.800 56.200 15.200 ;
        RECT 55.000 12.200 55.300 14.800 ;
        RECT 55.000 11.800 55.400 12.200 ;
        RECT 47.000 8.800 47.400 9.200 ;
        RECT 48.600 9.100 48.900 11.800 ;
        RECT 50.200 9.200 50.500 11.800 ;
        RECT 48.600 8.800 49.700 9.100 ;
        RECT 50.200 8.800 50.600 9.200 ;
        RECT 46.200 7.100 46.600 7.200 ;
        RECT 47.000 7.100 47.300 8.800 ;
        RECT 49.400 8.200 49.700 8.800 ;
        RECT 46.200 6.800 47.300 7.100 ;
        RECT 48.600 7.800 49.000 8.200 ;
        RECT 49.400 7.800 49.800 8.200 ;
        RECT 51.800 7.800 52.200 8.200 ;
        RECT 45.400 5.800 45.800 6.200 ;
        RECT 48.600 5.200 48.900 7.800 ;
        RECT 51.800 7.200 52.100 7.800 ;
        RECT 51.800 6.800 52.200 7.200 ;
        RECT 49.400 5.800 49.800 6.200 ;
        RECT 51.000 5.800 51.400 6.200 ;
        RECT 53.400 5.800 53.800 6.200 ;
        RECT 49.400 5.200 49.700 5.800 ;
        RECT 51.000 5.200 51.300 5.800 ;
        RECT 48.600 4.800 49.000 5.200 ;
        RECT 49.400 4.800 49.800 5.200 ;
        RECT 51.000 4.800 51.400 5.200 ;
        RECT 53.400 4.200 53.700 5.800 ;
        RECT 55.800 5.200 56.100 14.800 ;
        RECT 56.600 12.100 57.000 17.900 ;
        RECT 57.400 13.800 57.800 14.200 ;
        RECT 57.400 13.200 57.700 13.800 ;
        RECT 57.400 12.800 57.800 13.200 ;
        RECT 58.200 13.100 58.600 15.900 ;
        RECT 59.800 15.800 60.200 16.200 ;
        RECT 59.800 14.200 60.100 15.800 ;
        RECT 59.000 14.100 59.400 14.200 ;
        RECT 59.800 14.100 60.200 14.200 ;
        RECT 59.000 13.800 60.200 14.100 ;
        RECT 61.400 12.800 61.800 13.200 ;
        RECT 60.600 8.800 61.000 9.200 ;
        RECT 60.600 8.200 60.900 8.800 ;
        RECT 61.400 8.200 61.700 12.800 ;
        RECT 62.200 10.200 62.500 31.800 ;
        RECT 66.200 30.100 66.500 32.800 ;
        RECT 65.400 29.800 66.500 30.100 ;
        RECT 63.000 25.100 63.400 27.900 ;
        RECT 65.400 26.200 65.700 29.800 ;
        RECT 69.400 27.800 69.800 28.200 ;
        RECT 71.800 27.800 72.200 28.200 ;
        RECT 65.400 25.800 65.800 26.200 ;
        RECT 69.400 25.200 69.700 27.800 ;
        RECT 71.800 26.200 72.100 27.800 ;
        RECT 75.000 26.200 75.300 33.800 ;
        RECT 78.200 33.100 78.600 33.200 ;
        RECT 79.000 33.100 79.400 33.200 ;
        RECT 79.800 33.100 80.200 35.900 ;
        RECT 78.200 32.800 79.400 33.100 ;
        RECT 71.800 25.800 72.200 26.200 ;
        RECT 74.200 26.100 74.600 26.200 ;
        RECT 75.000 26.100 75.400 26.200 ;
        RECT 74.200 25.800 75.400 26.100 ;
        RECT 76.600 26.100 77.000 26.200 ;
        RECT 77.400 26.100 77.800 26.200 ;
        RECT 76.600 25.800 77.800 26.100 ;
        RECT 69.400 24.800 69.800 25.200 ;
        RECT 71.800 23.200 72.100 25.800 ;
        RECT 73.400 24.800 73.800 25.200 ;
        RECT 73.400 24.200 73.700 24.800 ;
        RECT 78.200 24.200 78.500 32.800 ;
        RECT 81.400 32.100 81.800 37.900 ;
        RECT 83.800 34.200 84.100 52.800 ;
        RECT 85.400 51.800 85.800 52.200 ;
        RECT 84.600 44.800 85.000 45.200 ;
        RECT 84.600 44.200 84.900 44.800 ;
        RECT 84.600 43.800 85.000 44.200 ;
        RECT 85.400 35.200 85.700 51.800 ;
        RECT 86.200 49.200 86.500 52.800 ;
        RECT 88.600 49.800 89.000 50.200 ;
        RECT 88.600 49.200 88.900 49.800 ;
        RECT 86.200 48.800 86.600 49.200 ;
        RECT 88.600 48.800 89.000 49.200 ;
        RECT 90.200 48.200 90.500 52.800 ;
        RECT 90.200 47.800 90.600 48.200 ;
        RECT 91.800 47.200 92.100 52.800 ;
        RECT 93.400 49.200 93.700 52.800 ;
        RECT 93.400 48.800 93.800 49.200 ;
        RECT 87.800 46.800 88.200 47.200 ;
        RECT 90.200 46.800 90.600 47.200 ;
        RECT 91.800 46.800 92.200 47.200 ;
        RECT 92.600 46.800 93.000 47.200 ;
        RECT 87.800 39.100 88.100 46.800 ;
        RECT 90.200 46.200 90.500 46.800 ;
        RECT 90.200 45.800 90.600 46.200 ;
        RECT 91.800 45.200 92.100 46.800 ;
        RECT 92.600 46.200 92.900 46.800 ;
        RECT 95.000 46.200 95.300 52.800 ;
        RECT 92.600 45.800 93.000 46.200 ;
        RECT 95.000 45.800 95.400 46.200 ;
        RECT 90.200 45.100 90.600 45.200 ;
        RECT 91.000 45.100 91.400 45.200 ;
        RECT 90.200 44.800 91.400 45.100 ;
        RECT 91.800 44.800 92.200 45.200 ;
        RECT 88.600 39.100 89.000 39.200 ;
        RECT 87.800 38.800 89.000 39.100 ;
        RECT 84.600 35.100 85.000 35.200 ;
        RECT 85.400 35.100 85.800 35.200 ;
        RECT 84.600 34.800 85.800 35.100 ;
        RECT 83.800 33.800 84.200 34.200 ;
        RECT 73.400 23.800 73.800 24.200 ;
        RECT 74.200 23.800 74.600 24.200 ;
        RECT 75.000 24.100 75.400 24.200 ;
        RECT 75.800 24.100 76.200 24.200 ;
        RECT 75.000 23.800 76.200 24.100 ;
        RECT 78.200 23.800 78.600 24.200 ;
        RECT 74.200 23.200 74.500 23.800 ;
        RECT 71.800 22.800 72.200 23.200 ;
        RECT 74.200 22.800 74.600 23.200 ;
        RECT 80.600 23.100 81.000 28.900 ;
        RECT 83.800 27.200 84.100 33.800 ;
        RECT 86.200 32.100 86.600 37.900 ;
        RECT 89.400 33.100 89.800 35.900 ;
        RECT 91.000 32.100 91.400 37.900 ;
        RECT 91.800 35.800 92.200 36.200 ;
        RECT 91.800 35.100 92.100 35.800 ;
        RECT 91.800 34.700 92.200 35.100 ;
        RECT 95.000 33.200 95.300 45.800 ;
        RECT 95.800 39.200 96.100 53.800 ;
        RECT 103.000 53.200 103.300 53.800 ;
        RECT 103.000 52.800 103.400 53.200 ;
        RECT 97.400 52.100 97.800 52.200 ;
        RECT 98.200 52.100 98.600 52.200 ;
        RECT 97.400 51.800 98.600 52.100 ;
        RECT 101.400 51.800 101.800 52.200 ;
        RECT 99.800 49.100 100.200 49.200 ;
        RECT 100.600 49.100 101.000 49.200 ;
        RECT 99.800 48.800 101.000 49.100 ;
        RECT 99.800 47.800 100.200 48.200 ;
        RECT 99.000 45.800 99.400 46.200 ;
        RECT 99.000 45.200 99.300 45.800 ;
        RECT 99.000 44.800 99.400 45.200 ;
        RECT 99.800 39.200 100.100 47.800 ;
        RECT 101.400 46.200 101.700 51.800 ;
        RECT 106.200 48.200 106.500 54.800 ;
        RECT 109.400 54.200 109.700 54.800 ;
        RECT 108.600 53.800 109.000 54.200 ;
        RECT 109.400 53.800 109.800 54.200 ;
        RECT 107.800 52.800 108.200 53.200 ;
        RECT 103.000 47.800 103.400 48.200 ;
        RECT 106.200 48.100 106.600 48.200 ;
        RECT 107.000 48.100 107.400 48.200 ;
        RECT 106.200 47.800 107.400 48.100 ;
        RECT 103.000 46.200 103.300 47.800 ;
        RECT 107.800 47.200 108.100 52.800 ;
        RECT 104.600 46.800 105.000 47.200 ;
        RECT 107.000 47.100 107.400 47.200 ;
        RECT 107.800 47.100 108.200 47.200 ;
        RECT 107.000 46.800 108.200 47.100 ;
        RECT 101.400 45.800 101.800 46.200 ;
        RECT 103.000 45.800 103.400 46.200 ;
        RECT 95.800 38.800 96.200 39.200 ;
        RECT 97.400 39.100 97.800 39.200 ;
        RECT 98.200 39.100 98.600 39.200 ;
        RECT 97.400 38.800 98.600 39.100 ;
        RECT 99.800 38.800 100.200 39.200 ;
        RECT 91.800 32.800 92.200 33.200 ;
        RECT 95.000 32.800 95.400 33.200 ;
        RECT 83.800 26.800 84.200 27.200 ;
        RECT 84.600 25.900 85.000 26.300 ;
        RECT 81.400 23.800 81.800 24.200 ;
        RECT 78.200 22.100 78.600 22.200 ;
        RECT 79.000 22.100 79.400 22.200 ;
        RECT 78.200 21.800 79.400 22.100 ;
        RECT 80.600 21.800 81.000 22.200 ;
        RECT 66.200 13.100 66.600 15.900 ;
        RECT 67.000 15.800 67.400 16.200 ;
        RECT 67.000 14.200 67.300 15.800 ;
        RECT 67.000 13.800 67.400 14.200 ;
        RECT 67.800 12.100 68.200 17.900 ;
        RECT 69.400 16.800 69.800 17.200 ;
        RECT 69.400 15.200 69.700 16.800 ;
        RECT 69.400 14.800 69.800 15.200 ;
        RECT 63.800 10.800 64.200 11.200 ;
        RECT 62.200 9.800 62.600 10.200 ;
        RECT 63.800 9.200 64.100 10.800 ;
        RECT 67.000 9.800 67.400 10.200 ;
        RECT 63.800 8.800 64.200 9.200 ;
        RECT 60.600 7.800 61.000 8.200 ;
        RECT 61.400 7.800 61.800 8.200 ;
        RECT 59.000 6.800 59.400 7.200 ;
        RECT 59.800 6.800 60.200 7.200 ;
        RECT 61.400 7.100 61.800 7.200 ;
        RECT 62.200 7.100 62.600 7.200 ;
        RECT 61.400 6.800 62.600 7.100 ;
        RECT 59.000 6.200 59.300 6.800 ;
        RECT 59.800 6.200 60.100 6.800 ;
        RECT 59.000 5.800 59.400 6.200 ;
        RECT 59.800 5.800 60.200 6.200 ;
        RECT 63.800 5.800 64.200 6.200 ;
        RECT 63.800 5.200 64.100 5.800 ;
        RECT 54.200 5.100 54.600 5.200 ;
        RECT 55.000 5.100 55.400 5.200 ;
        RECT 54.200 4.800 55.400 5.100 ;
        RECT 55.800 4.800 56.200 5.200 ;
        RECT 63.800 4.800 64.200 5.200 ;
        RECT 64.600 5.100 65.000 7.900 ;
        RECT 53.400 3.800 53.800 4.200 ;
        RECT 66.200 3.100 66.600 8.900 ;
        RECT 67.000 8.200 67.300 9.800 ;
        RECT 67.000 7.800 67.400 8.200 ;
        RECT 69.400 6.200 69.700 14.800 ;
        RECT 72.600 12.100 73.000 17.900 ;
        RECT 75.800 17.800 76.200 18.200 ;
        RECT 75.800 17.200 76.100 17.800 ;
        RECT 75.800 16.800 76.200 17.200 ;
        RECT 75.000 15.800 75.400 16.200 ;
        RECT 77.400 16.100 77.800 16.200 ;
        RECT 78.200 16.100 78.600 16.200 ;
        RECT 77.400 15.800 78.600 16.100 ;
        RECT 75.000 12.200 75.300 15.800 ;
        RECT 77.400 14.800 77.800 15.200 ;
        RECT 75.000 12.100 75.400 12.200 ;
        RECT 74.200 11.800 75.400 12.100 ;
        RECT 69.400 5.800 69.800 6.200 ;
        RECT 71.000 3.100 71.400 8.900 ;
        RECT 74.200 8.200 74.500 11.800 ;
        RECT 77.400 9.200 77.700 14.800 ;
        RECT 80.600 14.200 80.900 21.800 ;
        RECT 81.400 19.200 81.700 23.800 ;
        RECT 84.600 19.200 84.900 25.900 ;
        RECT 85.400 23.100 85.800 28.900 ;
        RECT 87.000 25.100 87.400 27.900 ;
        RECT 90.200 23.100 90.600 28.900 ;
        RECT 91.800 27.200 92.100 32.800 ;
        RECT 95.800 32.100 96.200 37.900 ;
        RECT 101.400 34.300 101.800 34.400 ;
        RECT 102.200 34.300 102.600 34.400 ;
        RECT 99.000 33.800 99.400 34.200 ;
        RECT 101.400 34.000 102.600 34.300 ;
        RECT 104.600 34.200 104.900 46.800 ;
        RECT 108.600 46.200 108.900 53.800 ;
        RECT 108.600 45.800 109.000 46.200 ;
        RECT 110.200 44.200 110.500 56.800 ;
        RECT 115.800 56.200 116.100 56.800 ;
        RECT 111.800 55.800 112.200 56.200 ;
        RECT 115.800 55.800 116.200 56.200 ;
        RECT 111.800 55.200 112.100 55.800 ;
        RECT 111.800 54.800 112.200 55.200 ;
        RECT 112.600 54.800 113.000 55.200 ;
        RECT 113.400 55.100 113.800 55.200 ;
        RECT 114.200 55.100 114.600 55.200 ;
        RECT 113.400 54.800 114.600 55.100 ;
        RECT 117.400 54.800 117.800 55.200 ;
        RECT 119.000 55.100 119.400 55.200 ;
        RECT 121.400 55.100 121.800 55.200 ;
        RECT 122.200 55.100 122.600 55.200 ;
        RECT 119.000 54.800 120.100 55.100 ;
        RECT 121.400 54.800 122.600 55.100 ;
        RECT 112.600 54.200 112.900 54.800 ;
        RECT 117.400 54.200 117.700 54.800 ;
        RECT 119.800 54.200 120.100 54.800 ;
        RECT 112.600 53.800 113.000 54.200 ;
        RECT 114.200 54.100 114.600 54.200 ;
        RECT 113.400 53.800 114.600 54.100 ;
        RECT 117.400 53.800 117.800 54.200 ;
        RECT 118.200 53.800 118.600 54.200 ;
        RECT 119.000 53.800 119.400 54.200 ;
        RECT 119.800 53.800 120.200 54.200 ;
        RECT 120.600 54.100 121.000 54.200 ;
        RECT 121.400 54.100 121.800 54.200 ;
        RECT 120.600 53.800 121.800 54.100 ;
        RECT 113.400 53.200 113.700 53.800 ;
        RECT 118.200 53.200 118.500 53.800 ;
        RECT 113.400 52.800 113.800 53.200 ;
        RECT 115.000 52.800 115.400 53.200 ;
        RECT 118.200 52.800 118.600 53.200 ;
        RECT 111.800 50.800 112.200 51.200 ;
        RECT 111.800 49.200 112.100 50.800 ;
        RECT 111.800 48.800 112.200 49.200 ;
        RECT 113.400 47.200 113.700 52.800 ;
        RECT 114.200 51.800 114.600 52.200 ;
        RECT 113.400 46.800 113.800 47.200 ;
        RECT 110.200 43.800 110.600 44.200 ;
        RECT 106.200 38.800 106.600 39.200 ;
        RECT 106.200 35.200 106.500 38.800 ;
        RECT 110.200 35.200 110.500 43.800 ;
        RECT 111.800 36.800 112.200 37.200 ;
        RECT 112.600 36.800 113.000 37.200 ;
        RECT 106.200 34.800 106.600 35.200 ;
        RECT 110.200 34.800 110.600 35.200 ;
        RECT 103.000 34.100 103.400 34.200 ;
        RECT 103.800 34.100 104.200 34.200 ;
        RECT 103.000 33.800 104.200 34.100 ;
        RECT 104.600 33.800 105.000 34.200 ;
        RECT 105.400 33.800 105.800 34.200 ;
        RECT 91.800 26.800 92.200 27.200 ;
        RECT 93.400 25.800 93.800 26.200 ;
        RECT 87.000 22.100 87.400 22.200 ;
        RECT 87.800 22.100 88.200 22.200 ;
        RECT 87.000 21.800 88.200 22.100 ;
        RECT 91.800 21.800 92.200 22.200 ;
        RECT 91.800 19.200 92.100 21.800 ;
        RECT 93.400 19.200 93.700 25.800 ;
        RECT 95.000 23.100 95.400 28.900 ;
        RECT 95.800 27.800 96.200 28.200 ;
        RECT 95.800 27.200 96.100 27.800 ;
        RECT 95.800 26.800 96.200 27.200 ;
        RECT 96.600 25.100 97.000 27.900 ;
        RECT 99.000 27.200 99.300 33.800 ;
        RECT 103.800 33.100 104.200 33.200 ;
        RECT 104.600 33.100 105.000 33.200 ;
        RECT 103.800 32.800 105.000 33.100 ;
        RECT 105.400 32.200 105.700 33.800 ;
        RECT 111.800 33.200 112.100 36.800 ;
        RECT 112.600 33.200 112.900 36.800 ;
        RECT 113.400 34.200 113.700 46.800 ;
        RECT 114.200 36.200 114.500 51.800 ;
        RECT 115.000 49.200 115.300 52.800 ;
        RECT 119.000 52.100 119.300 53.800 ;
        RECT 118.200 51.800 119.300 52.100 ;
        RECT 118.200 49.200 118.500 51.800 ;
        RECT 115.000 48.800 115.400 49.200 ;
        RECT 118.200 48.800 118.600 49.200 ;
        RECT 119.000 48.800 119.400 49.200 ;
        RECT 119.800 48.800 120.200 49.200 ;
        RECT 119.000 48.200 119.300 48.800 ;
        RECT 119.000 47.800 119.400 48.200 ;
        RECT 119.800 47.200 120.100 48.800 ;
        RECT 119.800 46.800 120.200 47.200 ;
        RECT 115.000 46.100 115.400 46.200 ;
        RECT 115.800 46.100 116.200 46.200 ;
        RECT 115.000 45.800 116.200 46.100 ;
        RECT 115.800 45.200 116.100 45.800 ;
        RECT 115.800 44.800 116.200 45.200 ;
        RECT 114.200 35.800 114.600 36.200 ;
        RECT 113.400 33.800 113.800 34.200 ;
        RECT 110.200 32.800 110.600 33.200 ;
        RECT 111.800 32.800 112.200 33.200 ;
        RECT 112.600 32.800 113.000 33.200 ;
        RECT 105.400 31.800 105.800 32.200 ;
        RECT 108.600 30.800 109.000 31.200 ;
        RECT 99.000 26.800 99.400 27.200 ;
        RECT 104.600 23.100 105.000 28.900 ;
        RECT 108.600 28.200 108.900 30.800 ;
        RECT 105.400 27.800 105.800 28.200 ;
        RECT 108.600 27.800 109.000 28.200 ;
        RECT 105.400 27.200 105.700 27.800 ;
        RECT 105.400 26.800 105.800 27.200 ;
        RECT 108.600 25.900 109.000 26.300 ;
        RECT 102.200 21.800 102.600 22.200 ;
        RECT 102.200 21.200 102.500 21.800 ;
        RECT 102.200 20.800 102.600 21.200 ;
        RECT 108.600 20.200 108.900 25.900 ;
        RECT 109.400 23.100 109.800 28.900 ;
        RECT 108.600 19.800 109.000 20.200 ;
        RECT 81.400 18.800 81.800 19.200 ;
        RECT 84.600 18.800 85.000 19.200 ;
        RECT 87.800 18.800 88.200 19.200 ;
        RECT 91.800 18.800 92.200 19.200 ;
        RECT 93.400 18.800 93.800 19.200 ;
        RECT 87.800 18.200 88.100 18.800 ;
        RECT 87.800 17.800 88.200 18.200 ;
        RECT 81.400 15.800 81.800 16.200 ;
        RECT 88.600 15.800 89.000 16.200 ;
        RECT 106.200 15.800 106.600 16.200 ;
        RECT 109.400 15.800 109.800 16.200 ;
        RECT 81.400 15.200 81.700 15.800 ;
        RECT 88.600 15.200 88.900 15.800 ;
        RECT 81.400 14.800 81.800 15.200 ;
        RECT 88.600 14.800 89.000 15.200 ;
        RECT 90.200 14.800 90.600 15.200 ;
        RECT 91.800 14.800 92.200 15.200 ;
        RECT 100.600 14.800 101.000 15.200 ;
        RECT 79.000 13.800 79.400 14.200 ;
        RECT 80.600 14.100 81.000 14.200 ;
        RECT 81.400 14.100 81.800 14.200 ;
        RECT 80.600 13.800 81.800 14.100 ;
        RECT 83.800 13.800 84.200 14.200 ;
        RECT 86.200 13.800 86.600 14.200 ;
        RECT 87.000 13.800 87.400 14.200 ;
        RECT 78.200 12.800 78.600 13.200 ;
        RECT 75.000 8.800 75.400 9.200 ;
        RECT 77.400 8.800 77.800 9.200 ;
        RECT 75.000 8.200 75.300 8.800 ;
        RECT 78.200 8.200 78.500 12.800 ;
        RECT 79.000 12.200 79.300 13.800 ;
        RECT 83.800 13.200 84.100 13.800 ;
        RECT 79.800 12.800 80.200 13.200 ;
        RECT 82.200 13.100 82.600 13.200 ;
        RECT 83.000 13.100 83.400 13.200 ;
        RECT 82.200 12.800 83.400 13.100 ;
        RECT 83.800 12.800 84.200 13.200 ;
        RECT 79.000 11.800 79.400 12.200 ;
        RECT 79.800 11.200 80.100 12.800 ;
        RECT 81.400 11.800 81.800 12.200 ;
        RECT 82.200 11.800 82.600 12.200 ;
        RECT 79.800 10.800 80.200 11.200 ;
        RECT 81.400 10.200 81.700 11.800 ;
        RECT 82.200 11.200 82.500 11.800 ;
        RECT 82.200 10.800 82.600 11.200 ;
        RECT 81.400 9.800 81.800 10.200 ;
        RECT 81.400 9.200 81.700 9.800 ;
        RECT 79.000 8.800 79.400 9.200 ;
        RECT 81.400 8.800 81.800 9.200 ;
        RECT 79.000 8.200 79.300 8.800 ;
        RECT 82.200 8.200 82.500 10.800 ;
        RECT 86.200 10.200 86.500 13.800 ;
        RECT 86.200 9.800 86.600 10.200 ;
        RECT 87.000 9.200 87.300 13.800 ;
        RECT 90.200 12.200 90.500 14.800 ;
        RECT 91.800 14.200 92.100 14.800 ;
        RECT 100.600 14.200 100.900 14.800 ;
        RECT 91.000 14.100 91.400 14.200 ;
        RECT 91.800 14.100 92.200 14.200 ;
        RECT 91.000 13.800 92.200 14.100 ;
        RECT 99.000 13.800 99.400 14.200 ;
        RECT 100.600 13.800 101.000 14.200 ;
        RECT 103.800 13.800 104.200 14.200 ;
        RECT 92.600 13.100 93.000 13.200 ;
        RECT 93.400 13.100 93.800 13.200 ;
        RECT 92.600 12.800 93.800 13.100 ;
        RECT 99.000 12.200 99.300 13.800 ;
        RECT 100.600 12.800 101.000 13.200 ;
        RECT 100.600 12.200 100.900 12.800 ;
        RECT 90.200 11.800 90.600 12.200 ;
        RECT 99.000 11.800 99.400 12.200 ;
        RECT 99.800 11.800 100.200 12.200 ;
        RECT 100.600 11.800 101.000 12.200 ;
        RECT 86.200 9.100 86.600 9.200 ;
        RECT 87.000 9.100 87.400 9.200 ;
        RECT 86.200 8.800 87.400 9.100 ;
        RECT 74.200 7.800 74.600 8.200 ;
        RECT 75.000 7.800 75.400 8.200 ;
        RECT 78.200 7.800 78.600 8.200 ;
        RECT 79.000 7.800 79.400 8.200 ;
        RECT 79.800 7.800 80.200 8.200 ;
        RECT 82.200 7.800 82.600 8.200 ;
        RECT 79.000 7.200 79.300 7.800 ;
        RECT 79.800 7.200 80.100 7.800 ;
        RECT 76.600 7.100 77.000 7.200 ;
        RECT 77.400 7.100 77.800 7.200 ;
        RECT 76.600 6.800 77.800 7.100 ;
        RECT 79.000 6.800 79.400 7.200 ;
        RECT 79.800 6.800 80.200 7.200 ;
        RECT 85.400 6.800 85.800 7.200 ;
        RECT 87.800 7.100 88.200 7.200 ;
        RECT 88.600 7.100 89.000 7.200 ;
        RECT 87.800 6.800 89.000 7.100 ;
        RECT 85.400 6.200 85.700 6.800 ;
        RECT 85.400 5.800 85.800 6.200 ;
        RECT 85.400 4.800 85.800 5.200 ;
        RECT 87.000 5.100 87.400 5.200 ;
        RECT 87.800 5.100 88.200 5.200 ;
        RECT 89.400 5.100 89.800 7.900 ;
        RECT 87.000 4.800 88.200 5.100 ;
        RECT 85.400 4.200 85.700 4.800 ;
        RECT 84.600 3.800 85.000 4.200 ;
        RECT 85.400 3.800 85.800 4.200 ;
        RECT 84.600 3.200 84.900 3.800 ;
        RECT 84.600 2.800 85.000 3.200 ;
        RECT 91.000 3.100 91.400 8.900 ;
        RECT 91.800 8.800 92.200 9.200 ;
        RECT 91.800 8.200 92.100 8.800 ;
        RECT 91.800 7.800 92.200 8.200 ;
        RECT 92.600 7.800 93.000 8.200 ;
        RECT 92.600 6.200 92.900 7.800 ;
        RECT 92.600 5.800 93.000 6.200 ;
        RECT 95.800 3.100 96.200 8.900 ;
        RECT 99.800 7.200 100.100 11.800 ;
        RECT 103.800 11.200 104.100 13.800 ;
        RECT 104.600 12.100 105.000 12.200 ;
        RECT 105.400 12.100 105.800 12.200 ;
        RECT 104.600 11.800 105.800 12.100 ;
        RECT 106.200 11.200 106.500 15.800 ;
        RECT 109.400 15.200 109.700 15.800 ;
        RECT 110.200 15.200 110.500 32.800 ;
        RECT 115.000 32.100 115.400 37.900 ;
        RECT 118.200 36.800 118.600 37.200 ;
        RECT 111.000 25.100 111.400 27.900 ;
        RECT 113.400 23.800 113.800 24.200 ;
        RECT 111.800 21.800 112.200 22.200 ;
        RECT 111.800 21.200 112.100 21.800 ;
        RECT 111.800 20.800 112.200 21.200 ;
        RECT 111.000 19.800 111.400 20.200 ;
        RECT 111.000 19.200 111.300 19.800 ;
        RECT 111.000 18.800 111.400 19.200 ;
        RECT 109.400 14.800 109.800 15.200 ;
        RECT 110.200 14.800 110.600 15.200 ;
        RECT 107.000 14.100 107.400 14.200 ;
        RECT 107.800 14.100 108.200 14.200 ;
        RECT 107.000 13.800 108.200 14.100 ;
        RECT 111.800 13.200 112.100 20.800 ;
        RECT 111.800 12.800 112.200 13.200 ;
        RECT 103.800 10.800 104.200 11.200 ;
        RECT 105.400 10.800 105.800 11.200 ;
        RECT 106.200 10.800 106.600 11.200 ;
        RECT 105.400 9.200 105.700 10.800 ;
        RECT 100.600 8.800 101.000 9.200 ;
        RECT 103.000 9.100 103.400 9.200 ;
        RECT 103.800 9.100 104.200 9.200 ;
        RECT 103.000 8.800 104.200 9.100 ;
        RECT 105.400 8.800 105.800 9.200 ;
        RECT 100.600 8.200 100.900 8.800 ;
        RECT 100.600 7.800 101.000 8.200 ;
        RECT 99.800 6.800 100.200 7.200 ;
        RECT 100.600 7.100 101.000 7.200 ;
        RECT 101.400 7.100 101.800 7.200 ;
        RECT 100.600 6.800 101.800 7.100 ;
        RECT 102.200 6.800 102.600 7.200 ;
        RECT 104.600 6.800 105.000 7.200 ;
        RECT 107.000 6.800 107.400 7.200 ;
        RECT 102.200 6.200 102.500 6.800 ;
        RECT 104.600 6.200 104.900 6.800 ;
        RECT 107.000 6.200 107.300 6.800 ;
        RECT 98.200 5.800 98.600 6.200 ;
        RECT 102.200 5.800 102.600 6.200 ;
        RECT 104.600 5.800 105.000 6.200 ;
        RECT 107.000 5.800 107.400 6.200 ;
        RECT 108.600 5.800 109.000 6.200 ;
        RECT 98.200 4.200 98.500 5.800 ;
        RECT 103.000 4.800 103.400 5.200 ;
        RECT 103.000 4.200 103.300 4.800 ;
        RECT 107.000 4.200 107.300 5.800 ;
        RECT 108.600 4.200 108.900 5.800 ;
        RECT 98.200 3.800 98.600 4.200 ;
        RECT 103.000 3.800 103.400 4.200 ;
        RECT 107.000 3.800 107.400 4.200 ;
        RECT 108.600 3.800 109.000 4.200 ;
        RECT 111.000 3.100 111.400 8.900 ;
        RECT 111.800 7.200 112.100 12.800 ;
        RECT 113.400 7.200 113.700 23.800 ;
        RECT 114.200 23.100 114.600 28.900 ;
        RECT 118.200 28.200 118.500 36.800 ;
        RECT 119.000 35.800 119.400 36.200 ;
        RECT 119.000 35.100 119.300 35.800 ;
        RECT 119.000 34.700 119.400 35.100 ;
        RECT 119.800 32.100 120.200 37.900 ;
        RECT 120.600 35.200 120.900 53.800 ;
        RECT 121.400 52.800 121.800 53.200 ;
        RECT 121.400 44.200 121.700 52.800 ;
        RECT 123.800 52.100 124.200 52.200 ;
        RECT 124.600 52.100 125.000 52.200 ;
        RECT 127.000 52.100 127.400 57.900 ;
        RECT 129.400 54.200 129.700 61.800 ;
        RECT 139.800 58.200 140.100 61.800 ;
        RECT 147.000 59.200 147.300 65.800 ;
        RECT 159.800 64.200 160.100 66.800 ;
        RECT 164.600 66.200 164.900 66.800 ;
        RECT 164.600 65.800 165.000 66.200 ;
        RECT 164.600 65.200 164.900 65.800 ;
        RECT 160.600 64.800 161.000 65.200 ;
        RECT 164.600 64.800 165.000 65.200 ;
        RECT 159.800 63.800 160.200 64.200 ;
        RECT 147.000 58.800 147.400 59.200 ;
        RECT 130.200 54.800 130.600 55.200 ;
        RECT 130.200 54.200 130.500 54.800 ;
        RECT 127.800 53.800 128.200 54.200 ;
        RECT 129.400 53.800 129.800 54.200 ;
        RECT 130.200 53.800 130.600 54.200 ;
        RECT 123.800 51.800 125.000 52.100 ;
        RECT 121.400 43.800 121.800 44.200 ;
        RECT 121.400 37.200 121.700 43.800 ;
        RECT 122.200 43.100 122.600 48.900 ;
        RECT 124.600 46.800 125.000 47.200 ;
        RECT 126.200 46.800 126.600 47.200 ;
        RECT 124.600 39.200 124.900 46.800 ;
        RECT 126.200 46.300 126.500 46.800 ;
        RECT 126.200 45.900 126.600 46.300 ;
        RECT 127.000 43.100 127.400 48.900 ;
        RECT 127.800 47.200 128.100 53.800 ;
        RECT 131.800 52.100 132.200 57.900 ;
        RECT 139.800 57.800 140.200 58.200 ;
        RECT 140.600 57.800 141.000 58.200 ;
        RECT 149.400 57.800 149.800 58.200 ;
        RECT 133.400 53.100 133.800 55.900 ;
        RECT 136.600 54.800 137.000 55.200 ;
        RECT 136.600 53.200 136.900 54.800 ;
        RECT 139.000 53.800 139.400 54.200 ;
        RECT 136.600 52.800 137.000 53.200 ;
        RECT 137.400 52.800 137.800 53.200 ;
        RECT 135.000 51.800 135.400 52.200 ;
        RECT 127.800 46.800 128.200 47.200 ;
        RECT 128.600 45.100 129.000 47.900 ;
        RECT 129.400 45.100 129.800 47.900 ;
        RECT 130.200 46.800 130.600 47.200 ;
        RECT 124.600 38.800 125.000 39.200 ;
        RECT 121.400 36.800 121.800 37.200 ;
        RECT 120.600 34.800 121.000 35.200 ;
        RECT 120.600 33.800 121.000 34.200 ;
        RECT 120.600 31.200 120.900 33.800 ;
        RECT 121.400 33.100 121.800 35.900 ;
        RECT 123.800 35.800 124.200 36.200 ;
        RECT 123.800 35.200 124.100 35.800 ;
        RECT 123.800 34.800 124.200 35.200 ;
        RECT 122.200 32.800 122.600 33.200 ;
        RECT 120.600 30.800 121.000 31.200 ;
        RECT 122.200 29.200 122.500 32.800 ;
        RECT 127.000 32.100 127.400 37.900 ;
        RECT 130.200 35.200 130.500 46.800 ;
        RECT 131.000 43.100 131.400 48.900 ;
        RECT 135.000 47.200 135.300 51.800 ;
        RECT 137.400 49.200 137.700 52.800 ;
        RECT 139.000 51.200 139.300 53.800 ;
        RECT 140.600 53.200 140.900 57.800 ;
        RECT 147.800 56.800 148.200 57.200 ;
        RECT 143.800 55.800 144.200 56.200 ;
        RECT 140.600 52.800 141.000 53.200 ;
        RECT 139.000 50.800 139.400 51.200 ;
        RECT 135.000 46.800 135.400 47.200 ;
        RECT 132.600 46.100 133.000 46.200 ;
        RECT 133.400 46.100 133.800 46.200 ;
        RECT 132.600 45.800 133.800 46.100 ;
        RECT 135.800 43.100 136.200 48.900 ;
        RECT 137.400 48.800 137.800 49.200 ;
        RECT 139.000 49.100 139.400 49.200 ;
        RECT 139.800 49.100 140.200 49.200 ;
        RECT 139.000 48.800 140.200 49.100 ;
        RECT 141.400 43.100 141.800 48.900 ;
        RECT 143.800 48.200 144.100 55.800 ;
        RECT 144.600 55.100 145.000 55.200 ;
        RECT 145.400 55.100 145.800 55.200 ;
        RECT 144.600 54.800 145.800 55.100 ;
        RECT 147.000 54.800 147.400 55.200 ;
        RECT 147.000 54.200 147.300 54.800 ;
        RECT 147.000 53.800 147.400 54.200 ;
        RECT 147.800 53.200 148.100 56.800 ;
        RECT 149.400 56.200 149.700 57.800 ;
        RECT 149.400 55.800 149.800 56.200 ;
        RECT 155.000 55.900 155.400 56.300 ;
        RECT 158.300 55.900 158.700 56.300 ;
        RECT 151.000 54.800 151.400 55.200 ;
        RECT 152.600 54.800 153.000 55.200 ;
        RECT 147.800 52.800 148.200 53.200 ;
        RECT 151.000 49.100 151.300 54.800 ;
        RECT 152.600 54.200 152.900 54.800 ;
        RECT 155.000 54.200 155.300 55.900 ;
        RECT 157.000 54.200 157.400 54.300 ;
        RECT 143.800 47.800 144.200 48.200 ;
        RECT 144.600 46.800 145.000 47.200 ;
        RECT 145.400 46.800 145.800 47.200 ;
        RECT 144.600 39.200 144.900 46.800 ;
        RECT 145.400 46.300 145.700 46.800 ;
        RECT 145.400 45.900 145.800 46.300 ;
        RECT 146.200 43.100 146.600 48.900 ;
        RECT 150.200 48.800 151.300 49.100 ;
        RECT 151.800 53.800 152.200 54.200 ;
        RECT 152.600 53.800 153.000 54.200 ;
        RECT 155.000 53.900 157.400 54.200 ;
        RECT 151.800 53.200 152.100 53.800 ;
        RECT 151.800 52.800 152.200 53.200 ;
        RECT 150.200 48.200 150.500 48.800 ;
        RECT 147.800 45.100 148.200 47.900 ;
        RECT 150.200 47.800 150.600 48.200 ;
        RECT 151.000 47.800 151.400 48.200 ;
        RECT 151.000 47.200 151.300 47.800 ;
        RECT 151.000 46.800 151.400 47.200 ;
        RECT 151.800 46.200 152.100 52.800 ;
        RECT 152.600 49.200 152.900 53.800 ;
        RECT 155.000 53.500 155.300 53.900 ;
        RECT 155.700 53.500 156.100 53.600 ;
        RECT 157.400 53.500 157.800 53.600 ;
        RECT 158.400 53.500 158.700 55.900 ;
        RECT 159.000 54.800 159.400 55.200 ;
        RECT 159.000 54.200 159.300 54.800 ;
        RECT 159.000 53.800 159.400 54.200 ;
        RECT 155.000 53.100 155.400 53.500 ;
        RECT 155.700 53.200 157.800 53.500 ;
        RECT 155.800 52.800 156.200 53.200 ;
        RECT 156.600 52.200 156.900 53.200 ;
        RECT 158.300 53.100 158.700 53.500 ;
        RECT 155.800 51.800 156.200 52.200 ;
        RECT 156.600 51.800 157.000 52.200 ;
        RECT 152.600 48.800 153.000 49.200 ;
        RECT 152.600 48.100 153.000 48.200 ;
        RECT 153.400 48.100 153.800 48.200 ;
        RECT 152.600 47.800 153.800 48.100 ;
        RECT 152.600 46.800 153.000 47.200 ;
        RECT 152.600 46.200 152.900 46.800 ;
        RECT 155.800 46.200 156.100 51.800 ;
        RECT 156.600 49.200 156.900 51.800 ;
        RECT 159.800 51.200 160.100 63.800 ;
        RECT 160.600 63.200 160.900 64.800 ;
        RECT 163.000 64.100 163.400 64.200 ;
        RECT 163.800 64.100 164.200 64.200 ;
        RECT 163.000 63.800 164.200 64.100 ;
        RECT 160.600 62.800 161.000 63.200 ;
        RECT 162.200 62.800 162.600 63.200 ;
        RECT 162.200 59.200 162.500 62.800 ;
        RECT 162.200 58.800 162.600 59.200 ;
        RECT 163.800 57.800 164.200 58.200 ;
        RECT 163.000 56.800 163.400 57.200 ;
        RECT 163.000 56.200 163.300 56.800 ;
        RECT 160.600 55.800 161.000 56.200 ;
        RECT 163.000 55.800 163.400 56.200 ;
        RECT 160.600 55.200 160.900 55.800 ;
        RECT 163.800 55.200 164.100 57.800 ;
        RECT 160.600 54.800 161.000 55.200 ;
        RECT 163.800 54.800 164.200 55.200 ;
        RECT 164.600 54.800 165.000 55.200 ;
        RECT 161.400 53.800 161.800 54.200 ;
        RECT 161.400 53.200 161.700 53.800 ;
        RECT 161.400 52.800 161.800 53.200 ;
        RECT 159.800 50.800 160.200 51.200 ;
        RECT 156.600 48.800 157.000 49.200 ;
        RECT 158.200 49.100 158.600 49.200 ;
        RECT 159.000 49.100 159.400 49.200 ;
        RECT 158.200 48.800 159.400 49.100 ;
        RECT 158.200 46.200 158.500 48.800 ;
        RECT 151.800 45.800 152.200 46.200 ;
        RECT 152.600 45.800 153.000 46.200 ;
        RECT 154.200 46.100 154.600 46.200 ;
        RECT 155.000 46.100 155.400 46.200 ;
        RECT 154.200 45.800 155.400 46.100 ;
        RECT 155.800 45.800 156.200 46.200 ;
        RECT 156.600 46.100 157.000 46.200 ;
        RECT 157.400 46.100 157.800 46.200 ;
        RECT 156.600 45.800 157.800 46.100 ;
        RECT 158.200 45.800 158.600 46.200 ;
        RECT 157.400 44.800 157.800 45.200 ;
        RECT 155.800 44.100 156.200 44.200 ;
        RECT 156.600 44.100 157.000 44.200 ;
        RECT 155.800 43.800 157.000 44.100 ;
        RECT 155.000 42.800 155.400 43.200 ;
        RECT 144.600 38.800 145.000 39.200 ;
        RECT 130.200 34.800 130.600 35.200 ;
        RECT 129.400 33.800 129.800 34.200 ;
        RECT 129.400 31.200 129.700 33.800 ;
        RECT 131.800 32.100 132.200 37.900 ;
        RECT 133.400 33.100 133.800 35.900 ;
        RECT 144.600 33.800 145.000 34.200 ;
        RECT 144.600 32.200 144.900 33.800 ;
        RECT 147.800 33.100 148.200 35.900 ;
        RECT 144.600 31.800 145.000 32.200 ;
        RECT 149.400 32.100 149.800 37.900 ;
        RECT 151.000 35.100 151.400 35.200 ;
        RECT 151.800 35.100 152.200 35.200 ;
        RECT 151.000 34.800 152.200 35.100 ;
        RECT 150.200 32.800 150.600 33.200 ;
        RECT 123.800 30.800 124.200 31.200 ;
        RECT 129.400 30.800 129.800 31.200 ;
        RECT 135.000 30.800 135.400 31.200 ;
        RECT 123.800 29.200 124.100 30.800 ;
        RECT 118.200 27.800 118.600 28.200 ;
        RECT 117.400 25.800 117.800 26.200 ;
        RECT 117.400 20.200 117.700 25.800 ;
        RECT 119.000 23.100 119.400 28.900 ;
        RECT 122.200 28.800 122.600 29.200 ;
        RECT 123.800 28.800 124.200 29.200 ;
        RECT 120.600 25.100 121.000 27.900 ;
        RECT 133.400 25.800 133.800 26.200 ;
        RECT 133.400 25.200 133.700 25.800 ;
        RECT 133.400 24.800 133.800 25.200 ;
        RECT 134.200 25.100 134.600 27.900 ;
        RECT 135.000 27.200 135.300 30.800 ;
        RECT 135.000 26.800 135.400 27.200 ;
        RECT 135.800 23.100 136.200 28.900 ;
        RECT 137.400 25.800 137.800 26.200 ;
        RECT 137.400 24.200 137.700 25.800 ;
        RECT 137.400 23.800 137.800 24.200 ;
        RECT 140.600 23.100 141.000 28.900 ;
        RECT 144.600 27.200 144.900 31.800 ;
        RECT 144.600 26.800 145.000 27.200 ;
        RECT 145.400 25.100 145.800 27.900 ;
        RECT 141.400 23.800 141.800 24.200 ;
        RECT 145.400 23.800 145.800 24.200 ;
        RECT 123.800 21.800 124.200 22.200 ;
        RECT 117.400 19.800 117.800 20.200 ;
        RECT 123.800 19.100 124.100 21.800 ;
        RECT 123.800 18.800 124.900 19.100 ;
        RECT 115.000 14.800 115.400 15.200 ;
        RECT 117.400 15.100 117.800 15.200 ;
        RECT 117.400 14.800 118.500 15.100 ;
        RECT 115.000 11.200 115.300 14.800 ;
        RECT 115.800 11.800 116.200 12.200 ;
        RECT 115.000 10.800 115.400 11.200 ;
        RECT 115.800 10.200 116.100 11.800 ;
        RECT 115.800 9.800 116.200 10.200 ;
        RECT 118.200 9.200 118.500 14.800 ;
        RECT 119.000 14.800 119.400 15.200 ;
        RECT 119.000 14.200 119.300 14.800 ;
        RECT 119.000 13.800 119.400 14.200 ;
        RECT 123.000 12.800 123.400 13.200 ;
        RECT 120.600 11.800 121.000 12.200 ;
        RECT 120.600 10.200 120.900 11.800 ;
        RECT 120.600 9.800 121.000 10.200 ;
        RECT 115.000 7.800 115.400 8.200 ;
        RECT 111.800 6.800 112.200 7.200 ;
        RECT 113.400 6.800 113.800 7.200 ;
        RECT 115.000 6.300 115.300 7.800 ;
        RECT 115.000 5.900 115.400 6.300 ;
        RECT 115.800 3.100 116.200 8.900 ;
        RECT 118.200 8.800 118.600 9.200 ;
        RECT 117.400 5.100 117.800 7.900 ;
        RECT 119.800 6.800 120.200 7.200 ;
        RECT 119.800 6.200 120.100 6.800 ;
        RECT 120.600 6.200 120.900 9.800 ;
        RECT 123.000 9.200 123.300 12.800 ;
        RECT 123.800 12.100 124.200 17.900 ;
        RECT 124.600 15.200 124.900 18.800 ;
        RECT 127.800 15.800 128.200 16.200 ;
        RECT 124.600 14.800 125.000 15.200 ;
        RECT 125.400 14.800 125.800 15.200 ;
        RECT 127.800 15.100 128.100 15.800 ;
        RECT 121.400 8.800 121.800 9.200 ;
        RECT 123.000 8.800 123.400 9.200 ;
        RECT 121.400 8.200 121.700 8.800 ;
        RECT 121.400 7.800 121.800 8.200 ;
        RECT 122.200 8.100 122.600 8.200 ;
        RECT 123.000 8.100 123.400 8.200 ;
        RECT 122.200 7.800 123.400 8.100 ;
        RECT 124.600 7.800 125.000 8.200 ;
        RECT 124.600 7.200 124.900 7.800 ;
        RECT 122.200 6.800 122.600 7.200 ;
        RECT 124.600 6.800 125.000 7.200 ;
        RECT 118.200 5.800 118.600 6.200 ;
        RECT 119.800 5.800 120.200 6.200 ;
        RECT 120.600 5.800 121.000 6.200 ;
        RECT 118.200 5.200 118.500 5.800 ;
        RECT 122.200 5.200 122.500 6.800 ;
        RECT 123.000 5.800 123.400 6.200 ;
        RECT 123.000 5.200 123.300 5.800 ;
        RECT 125.400 5.200 125.700 14.800 ;
        RECT 127.800 14.700 128.200 15.100 ;
        RECT 128.600 12.100 129.000 17.900 ;
        RECT 133.400 16.100 133.800 16.200 ;
        RECT 134.200 16.100 134.600 16.200 ;
        RECT 130.200 13.100 130.600 15.900 ;
        RECT 133.400 15.800 134.600 16.100 ;
        RECT 139.000 16.100 139.400 16.200 ;
        RECT 139.800 16.100 140.200 16.200 ;
        RECT 139.000 15.800 140.200 16.100 ;
        RECT 131.800 14.800 132.200 15.200 ;
        RECT 131.000 13.800 131.400 14.200 ;
        RECT 131.000 13.200 131.300 13.800 ;
        RECT 131.000 12.800 131.400 13.200 ;
        RECT 131.800 12.200 132.100 14.800 ;
        RECT 131.800 11.800 132.200 12.200 ;
        RECT 126.200 8.800 126.600 9.200 ;
        RECT 126.200 7.200 126.500 8.800 ;
        RECT 126.200 6.800 126.600 7.200 ;
        RECT 126.200 6.100 126.600 6.200 ;
        RECT 127.000 6.100 127.400 6.200 ;
        RECT 126.200 5.800 127.400 6.100 ;
        RECT 127.800 5.800 128.200 6.200 ;
        RECT 127.800 5.200 128.100 5.800 ;
        RECT 118.200 4.800 118.600 5.200 ;
        RECT 122.200 4.800 122.600 5.200 ;
        RECT 123.000 4.800 123.400 5.200 ;
        RECT 125.400 5.100 125.800 5.200 ;
        RECT 126.200 5.100 126.600 5.200 ;
        RECT 125.400 4.800 126.600 5.100 ;
        RECT 127.800 4.800 128.200 5.200 ;
        RECT 128.600 5.100 129.000 7.900 ;
        RECT 129.400 7.800 129.800 8.200 ;
        RECT 129.400 7.200 129.700 7.800 ;
        RECT 129.400 6.800 129.800 7.200 ;
        RECT 130.200 3.100 130.600 8.900 ;
        RECT 131.800 6.200 132.100 11.800 ;
        RECT 131.800 5.800 132.200 6.200 ;
        RECT 133.400 5.200 133.700 15.800 ;
        RECT 141.400 15.200 141.700 23.800 ;
        RECT 143.000 21.800 143.400 22.200 ;
        RECT 143.000 19.200 143.300 21.800 ;
        RECT 143.000 18.800 143.400 19.200 ;
        RECT 135.000 14.800 135.400 15.200 ;
        RECT 136.600 14.800 137.000 15.200 ;
        RECT 137.400 14.800 137.800 15.200 ;
        RECT 139.000 14.800 139.400 15.200 ;
        RECT 139.800 14.800 140.200 15.200 ;
        RECT 141.400 14.800 141.800 15.200 ;
        RECT 135.000 10.200 135.300 14.800 ;
        RECT 136.600 14.200 136.900 14.800 ;
        RECT 135.800 13.800 136.200 14.200 ;
        RECT 136.600 13.800 137.000 14.200 ;
        RECT 135.800 12.200 136.100 13.800 ;
        RECT 135.800 11.800 136.200 12.200 ;
        RECT 137.400 10.200 137.700 14.800 ;
        RECT 139.000 14.200 139.300 14.800 ;
        RECT 139.000 13.800 139.400 14.200 ;
        RECT 139.800 11.200 140.100 14.800 ;
        RECT 140.600 13.800 141.000 14.200 ;
        RECT 142.200 13.800 142.600 14.200 ;
        RECT 140.600 12.200 140.900 13.800 ;
        RECT 142.200 13.200 142.500 13.800 ;
        RECT 142.200 12.800 142.600 13.200 ;
        RECT 143.000 13.100 143.400 15.900 ;
        RECT 143.800 14.800 144.200 15.200 ;
        RECT 140.600 11.800 141.000 12.200 ;
        RECT 141.400 11.800 141.800 12.200 ;
        RECT 139.800 10.800 140.200 11.200 ;
        RECT 135.000 9.800 135.400 10.200 ;
        RECT 137.400 9.800 137.800 10.200 ;
        RECT 139.000 9.800 139.400 10.200 ;
        RECT 136.600 9.100 137.000 9.200 ;
        RECT 137.400 9.100 137.800 9.200 ;
        RECT 133.400 4.800 133.800 5.200 ;
        RECT 135.000 3.100 135.400 8.900 ;
        RECT 136.600 8.800 137.800 9.100 ;
        RECT 139.000 6.200 139.300 9.800 ;
        RECT 139.800 9.100 140.100 10.800 ;
        RECT 141.400 9.200 141.700 11.800 ;
        RECT 140.600 9.100 141.000 9.200 ;
        RECT 139.800 8.800 141.000 9.100 ;
        RECT 141.400 8.800 141.800 9.200 ;
        RECT 139.000 5.800 139.400 6.200 ;
        RECT 141.400 5.100 141.800 7.900 ;
        RECT 143.000 3.100 143.400 8.900 ;
        RECT 143.800 8.200 144.100 14.800 ;
        RECT 144.600 12.100 145.000 17.900 ;
        RECT 145.400 15.100 145.700 23.800 ;
        RECT 147.000 23.100 147.400 28.900 ;
        RECT 148.600 26.100 149.000 26.200 ;
        RECT 149.400 26.100 149.800 26.200 ;
        RECT 148.600 25.800 149.800 26.100 ;
        RECT 148.600 22.200 148.900 25.800 ;
        RECT 148.600 21.800 149.000 22.200 ;
        RECT 145.400 14.700 145.800 15.100 ;
        RECT 145.400 12.800 145.800 13.200 ;
        RECT 144.600 8.800 145.000 9.200 ;
        RECT 143.800 7.800 144.200 8.200 ;
        RECT 144.600 6.200 144.900 8.800 ;
        RECT 145.400 8.200 145.700 12.800 ;
        RECT 149.400 12.100 149.800 17.900 ;
        RECT 150.200 17.200 150.500 32.800 ;
        RECT 154.200 32.100 154.600 37.900 ;
        RECT 155.000 29.200 155.300 42.800 ;
        RECT 156.600 39.200 156.900 43.800 ;
        RECT 157.400 43.200 157.700 44.800 ;
        RECT 159.800 43.800 160.200 44.200 ;
        RECT 157.400 42.800 157.800 43.200 ;
        RECT 156.600 38.800 157.000 39.200 ;
        RECT 157.400 33.100 157.800 35.900 ;
        RECT 158.200 33.800 158.600 34.200 ;
        RECT 158.200 33.200 158.500 33.800 ;
        RECT 158.200 32.800 158.600 33.200 ;
        RECT 154.200 29.100 154.600 29.200 ;
        RECT 155.000 29.100 155.400 29.200 ;
        RECT 151.800 23.100 152.200 28.900 ;
        RECT 154.200 28.800 155.400 29.100 ;
        RECT 155.000 25.100 155.400 27.900 ;
        RECT 156.600 23.100 157.000 28.900 ;
        RECT 157.400 25.900 157.800 26.300 ;
        RECT 157.400 25.200 157.700 25.900 ;
        RECT 157.400 24.800 157.800 25.200 ;
        RECT 151.800 19.100 152.200 19.200 ;
        RECT 152.600 19.100 153.000 19.200 ;
        RECT 151.800 18.800 153.000 19.100 ;
        RECT 150.200 16.800 150.600 17.200 ;
        RECT 154.200 15.800 154.600 16.200 ;
        RECT 154.200 14.200 154.500 15.800 ;
        RECT 155.000 15.100 155.400 15.200 ;
        RECT 155.800 15.100 156.200 15.200 ;
        RECT 155.000 14.800 156.200 15.100 ;
        RECT 158.200 14.200 158.500 32.800 ;
        RECT 159.000 32.100 159.400 37.900 ;
        RECT 159.800 26.200 160.100 43.800 ;
        RECT 160.600 43.100 161.000 48.900 ;
        RECT 161.400 44.200 161.700 52.800 ;
        RECT 162.200 49.800 162.600 50.200 ;
        RECT 161.400 43.800 161.800 44.200 ;
        RECT 162.200 35.200 162.500 49.800 ;
        RECT 164.600 49.200 164.900 54.800 ;
        RECT 165.400 53.800 165.800 54.200 ;
        RECT 165.400 52.200 165.700 53.800 ;
        RECT 165.400 51.800 165.800 52.200 ;
        RECT 164.600 48.800 165.000 49.200 ;
        RECT 163.800 46.200 164.200 46.300 ;
        RECT 164.600 46.200 165.000 46.300 ;
        RECT 163.800 45.900 165.000 46.200 ;
        RECT 165.400 43.100 165.800 48.900 ;
        RECT 166.200 47.200 166.500 66.800 ;
        RECT 170.200 66.200 170.500 66.800 ;
        RECT 170.200 65.800 170.600 66.200 ;
        RECT 169.400 64.800 169.800 65.200 ;
        RECT 169.400 64.200 169.700 64.800 ;
        RECT 169.400 63.800 169.800 64.200 ;
        RECT 171.800 62.800 172.200 63.200 ;
        RECT 167.000 61.800 167.400 62.200 ;
        RECT 167.000 58.200 167.300 61.800 ;
        RECT 167.000 57.800 167.400 58.200 ;
        RECT 170.200 57.800 170.600 58.200 ;
        RECT 171.000 57.800 171.400 58.200 ;
        RECT 170.200 56.200 170.500 57.800 ;
        RECT 171.000 56.200 171.300 57.800 ;
        RECT 171.800 57.200 172.100 62.800 ;
        RECT 171.800 56.800 172.200 57.200 ;
        RECT 171.800 56.200 172.100 56.800 ;
        RECT 167.000 55.800 167.400 56.200 ;
        RECT 169.400 55.800 169.800 56.200 ;
        RECT 170.200 55.800 170.600 56.200 ;
        RECT 171.000 55.800 171.400 56.200 ;
        RECT 171.800 55.800 172.200 56.200 ;
        RECT 167.000 55.200 167.300 55.800 ;
        RECT 169.400 55.200 169.700 55.800 ;
        RECT 167.000 54.800 167.400 55.200 ;
        RECT 169.400 54.800 169.800 55.200 ;
        RECT 171.000 54.800 171.400 55.200 ;
        RECT 171.000 54.200 171.300 54.800 ;
        RECT 172.600 54.200 172.900 73.800 ;
        RECT 173.400 73.200 173.700 76.800 ;
        RECT 174.200 75.200 174.500 81.800 ;
        RECT 178.200 77.200 178.500 81.800 ;
        RECT 178.200 76.800 178.600 77.200 ;
        RECT 174.200 74.800 174.600 75.200 ;
        RECT 173.400 72.800 173.800 73.200 ;
        RECT 175.800 73.100 176.200 73.200 ;
        RECT 176.600 73.100 177.000 73.200 ;
        RECT 175.800 72.800 177.000 73.100 ;
        RECT 177.400 72.800 177.800 73.200 ;
        RECT 173.400 70.200 173.700 72.800 ;
        RECT 175.800 71.800 176.200 72.200 ;
        RECT 173.400 69.800 173.800 70.200 ;
        RECT 173.400 68.200 173.700 69.800 ;
        RECT 173.400 67.800 173.800 68.200 ;
        RECT 175.800 67.100 176.100 71.800 ;
        RECT 177.400 71.200 177.700 72.800 ;
        RECT 178.200 71.800 178.600 72.200 ;
        RECT 177.400 70.800 177.800 71.200 ;
        RECT 176.600 67.100 177.000 67.200 ;
        RECT 175.800 66.800 177.000 67.100 ;
        RECT 178.200 66.200 178.500 71.800 ;
        RECT 179.000 69.200 179.300 85.800 ;
        RECT 182.200 85.100 182.500 86.800 ;
        RECT 184.200 86.700 184.600 86.800 ;
        RECT 182.200 84.700 182.600 85.100 ;
        RECT 183.800 84.800 184.200 85.200 ;
        RECT 185.600 85.100 185.900 87.500 ;
        RECT 180.600 76.800 181.000 77.200 ;
        RECT 180.600 76.200 180.900 76.800 ;
        RECT 179.800 75.800 180.200 76.200 ;
        RECT 180.600 75.800 181.000 76.200 ;
        RECT 179.800 75.200 180.100 75.800 ;
        RECT 179.800 74.800 180.200 75.200 ;
        RECT 183.800 73.200 184.100 84.800 ;
        RECT 185.500 84.700 185.900 85.100 ;
        RECT 186.200 86.800 186.600 87.200 ;
        RECT 186.200 83.200 186.500 86.800 ;
        RECT 191.800 86.200 192.100 90.800 ;
        RECT 191.800 85.800 192.200 86.200 ;
        RECT 186.200 82.800 186.600 83.200 ;
        RECT 183.800 72.800 184.200 73.200 ;
        RECT 184.600 73.100 185.000 75.900 ;
        RECT 185.400 74.800 185.800 75.200 ;
        RECT 185.400 74.200 185.700 74.800 ;
        RECT 185.400 73.800 185.800 74.200 ;
        RECT 183.800 69.200 184.100 72.800 ;
        RECT 186.200 72.100 186.600 77.900 ;
        RECT 187.000 74.700 187.400 75.100 ;
        RECT 179.000 68.800 179.400 69.200 ;
        RECT 179.000 68.200 179.300 68.800 ;
        RECT 179.000 67.800 179.400 68.200 ;
        RECT 173.400 66.100 173.800 66.200 ;
        RECT 174.200 66.100 174.600 66.200 ;
        RECT 173.400 65.800 174.600 66.100 ;
        RECT 175.000 66.100 175.400 66.200 ;
        RECT 175.800 66.100 176.200 66.200 ;
        RECT 175.000 65.800 176.200 66.100 ;
        RECT 176.600 65.800 177.000 66.200 ;
        RECT 178.200 65.800 178.600 66.200 ;
        RECT 173.400 65.100 173.800 65.200 ;
        RECT 174.200 65.100 174.600 65.200 ;
        RECT 173.400 64.800 174.600 65.100 ;
        RECT 175.800 65.100 176.200 65.200 ;
        RECT 176.600 65.100 176.900 65.800 ;
        RECT 179.800 65.100 180.200 67.900 ;
        RECT 180.600 67.800 181.000 68.200 ;
        RECT 180.600 67.200 180.900 67.800 ;
        RECT 180.600 66.800 181.000 67.200 ;
        RECT 175.800 64.800 176.900 65.100 ;
        RECT 181.400 63.100 181.800 68.900 ;
        RECT 183.800 68.800 184.200 69.200 ;
        RECT 182.200 66.800 182.600 67.200 ;
        RECT 182.200 66.300 182.500 66.800 ;
        RECT 182.200 65.900 182.600 66.300 ;
        RECT 186.200 63.100 186.600 68.900 ;
        RECT 187.000 67.200 187.300 74.700 ;
        RECT 191.000 72.100 191.400 77.900 ;
        RECT 193.400 71.800 193.800 72.200 ;
        RECT 192.600 69.800 193.000 70.200 ;
        RECT 187.800 69.100 188.200 69.200 ;
        RECT 188.600 69.100 189.000 69.200 ;
        RECT 187.800 68.800 189.000 69.100 ;
        RECT 187.000 66.800 187.400 67.200 ;
        RECT 187.000 63.800 187.400 64.200 ;
        RECT 178.200 61.800 178.600 62.200 ;
        RECT 178.200 57.200 178.500 61.800 ;
        RECT 178.200 56.800 178.600 57.200 ;
        RECT 179.800 56.100 180.200 56.200 ;
        RECT 180.600 56.100 181.000 56.200 ;
        RECT 179.800 55.800 181.000 56.100 ;
        RECT 175.000 55.100 175.400 55.200 ;
        RECT 175.800 55.100 176.200 55.200 ;
        RECT 175.000 54.800 176.200 55.100 ;
        RECT 176.600 55.100 177.000 55.200 ;
        RECT 177.400 55.100 177.800 55.200 ;
        RECT 176.600 54.800 177.800 55.100 ;
        RECT 179.800 54.800 180.200 55.200 ;
        RECT 182.200 54.800 182.600 55.200 ;
        RECT 167.800 53.800 168.200 54.200 ;
        RECT 171.000 53.800 171.400 54.200 ;
        RECT 172.600 53.800 173.000 54.200 ;
        RECT 176.600 54.100 177.000 54.200 ;
        RECT 177.400 54.100 177.800 54.200 ;
        RECT 176.600 53.800 177.800 54.100 ;
        RECT 178.200 54.100 178.600 54.200 ;
        RECT 179.000 54.100 179.400 54.200 ;
        RECT 178.200 53.800 179.400 54.100 ;
        RECT 166.200 46.800 166.600 47.200 ;
        RECT 167.000 45.100 167.400 47.900 ;
        RECT 167.800 45.200 168.100 53.800 ;
        RECT 172.600 53.100 173.000 53.200 ;
        RECT 173.400 53.100 173.800 53.200 ;
        RECT 172.600 52.800 173.800 53.100 ;
        RECT 178.200 52.800 178.600 53.200 ;
        RECT 168.600 51.800 169.000 52.200 ;
        RECT 168.600 50.200 168.900 51.800 ;
        RECT 168.600 49.800 169.000 50.200 ;
        RECT 171.800 49.800 172.200 50.200 ;
        RECT 168.600 48.100 169.000 48.200 ;
        RECT 169.400 48.100 169.800 48.200 ;
        RECT 170.200 48.100 170.600 48.200 ;
        RECT 168.600 47.800 170.600 48.100 ;
        RECT 168.600 47.100 169.000 47.200 ;
        RECT 169.400 47.100 169.800 47.200 ;
        RECT 168.600 46.800 169.800 47.100 ;
        RECT 171.800 46.200 172.100 49.800 ;
        RECT 170.200 46.100 170.600 46.200 ;
        RECT 171.000 46.100 171.400 46.200 ;
        RECT 170.200 45.800 171.400 46.100 ;
        RECT 171.800 45.800 172.200 46.200 ;
        RECT 167.800 45.100 168.200 45.200 ;
        RECT 168.600 45.100 169.000 45.200 ;
        RECT 172.600 45.100 173.000 47.900 ;
        RECT 173.400 46.800 173.800 47.200 ;
        RECT 167.800 44.800 169.000 45.100 ;
        RECT 166.200 43.800 166.600 44.200 ;
        RECT 166.200 39.200 166.500 43.800 ;
        RECT 166.200 38.800 166.600 39.200 ;
        RECT 162.200 34.800 162.600 35.200 ;
        RECT 163.800 32.100 164.200 37.900 ;
        RECT 167.800 35.100 168.200 35.200 ;
        RECT 168.600 35.100 169.000 35.200 ;
        RECT 167.800 34.800 169.000 35.100 ;
        RECT 168.600 33.800 169.000 34.200 ;
        RECT 167.000 32.800 167.400 33.200 ;
        RECT 167.000 29.200 167.300 32.800 ;
        RECT 167.800 29.800 168.200 30.200 ;
        RECT 167.800 29.200 168.100 29.800 ;
        RECT 159.800 25.800 160.200 26.200 ;
        RECT 154.200 14.100 154.600 14.200 ;
        RECT 155.000 14.100 155.400 14.200 ;
        RECT 154.200 13.800 155.400 14.100 ;
        RECT 157.400 13.800 157.800 14.200 ;
        RECT 158.200 13.800 158.600 14.200 ;
        RECT 154.200 13.100 154.600 13.200 ;
        RECT 155.000 13.100 155.400 13.200 ;
        RECT 154.200 12.800 155.400 13.100 ;
        RECT 150.200 9.800 150.600 10.200 ;
        RECT 150.200 9.200 150.500 9.800 ;
        RECT 145.400 7.800 145.800 8.200 ;
        RECT 144.600 5.800 145.000 6.200 ;
        RECT 147.800 3.100 148.200 8.900 ;
        RECT 150.200 8.800 150.600 9.200 ;
        RECT 155.000 3.100 155.400 8.900 ;
        RECT 157.400 6.200 157.700 13.800 ;
        RECT 158.200 12.800 158.600 13.200 ;
        RECT 159.000 13.100 159.400 15.900 ;
        RECT 158.200 12.200 158.500 12.800 ;
        RECT 158.200 11.800 158.600 12.200 ;
        RECT 159.800 10.100 160.100 25.800 ;
        RECT 161.400 23.100 161.800 28.900 ;
        RECT 162.200 28.800 162.600 29.200 ;
        RECT 164.600 29.100 165.000 29.200 ;
        RECT 165.400 29.100 165.800 29.200 ;
        RECT 164.600 28.800 165.800 29.100 ;
        RECT 167.000 28.800 167.400 29.200 ;
        RECT 167.800 28.800 168.200 29.200 ;
        RECT 162.200 28.200 162.500 28.800 ;
        RECT 168.600 28.200 168.900 33.800 ;
        RECT 170.200 31.800 170.600 32.200 ;
        RECT 172.600 32.100 173.000 37.900 ;
        RECT 173.400 35.200 173.700 46.800 ;
        RECT 174.200 43.100 174.600 48.900 ;
        RECT 175.000 46.800 175.400 47.200 ;
        RECT 175.000 46.300 175.300 46.800 ;
        RECT 175.000 45.900 175.400 46.300 ;
        RECT 178.200 43.200 178.500 52.800 ;
        RECT 178.200 42.800 178.600 43.200 ;
        RECT 179.000 43.100 179.400 48.900 ;
        RECT 179.800 46.200 180.100 54.800 ;
        RECT 182.200 54.200 182.500 54.800 ;
        RECT 182.200 53.800 182.600 54.200 ;
        RECT 183.000 53.800 183.400 54.200 ;
        RECT 180.600 51.800 181.000 52.200 ;
        RECT 180.600 50.200 180.900 51.800 ;
        RECT 180.600 49.800 181.000 50.200 ;
        RECT 180.600 49.100 181.000 49.200 ;
        RECT 181.400 49.100 181.800 49.200 ;
        RECT 180.600 48.800 181.800 49.100 ;
        RECT 179.800 45.800 180.200 46.200 ;
        RECT 182.200 45.100 182.600 47.900 ;
        RECT 173.400 34.800 173.800 35.200 ;
        RECT 174.200 34.800 174.600 35.200 ;
        RECT 175.000 35.100 175.400 35.200 ;
        RECT 175.800 35.100 176.200 35.200 ;
        RECT 175.000 34.800 176.200 35.100 ;
        RECT 173.400 34.200 173.700 34.800 ;
        RECT 173.400 33.800 173.800 34.200 ;
        RECT 170.200 30.200 170.500 31.800 ;
        RECT 170.200 29.800 170.600 30.200 ;
        RECT 162.200 27.800 162.600 28.200 ;
        RECT 167.000 27.800 167.400 28.200 ;
        RECT 168.600 27.800 169.000 28.200 ;
        RECT 167.000 27.200 167.300 27.800 ;
        RECT 167.000 26.800 167.400 27.200 ;
        RECT 168.600 26.800 169.000 27.200 ;
        RECT 164.600 24.800 165.000 25.200 ;
        RECT 160.600 12.100 161.000 17.900 ;
        RECT 163.000 14.800 163.400 15.200 ;
        RECT 159.000 9.800 160.100 10.100 ;
        RECT 162.200 11.800 162.600 12.200 ;
        RECT 158.200 8.800 158.600 9.200 ;
        RECT 158.200 6.200 158.500 8.800 ;
        RECT 159.000 8.200 159.300 9.800 ;
        RECT 162.200 9.200 162.500 11.800 ;
        RECT 159.000 7.800 159.400 8.200 ;
        RECT 159.000 7.200 159.300 7.800 ;
        RECT 159.000 6.800 159.400 7.200 ;
        RECT 157.400 5.800 157.800 6.200 ;
        RECT 158.200 5.800 158.600 6.200 ;
        RECT 159.800 3.100 160.200 8.900 ;
        RECT 162.200 8.800 162.600 9.200 ;
        RECT 162.200 8.200 162.500 8.800 ;
        RECT 163.000 8.200 163.300 14.800 ;
        RECT 164.600 14.200 164.900 24.800 ;
        RECT 164.600 13.800 165.000 14.200 ;
        RECT 165.400 12.100 165.800 17.900 ;
        RECT 168.600 16.200 168.900 26.800 ;
        RECT 170.200 23.100 170.600 28.900 ;
        RECT 174.200 26.300 174.500 34.800 ;
        RECT 177.400 32.100 177.800 37.900 ;
        RECT 179.000 33.100 179.400 35.900 ;
        RECT 179.800 33.100 180.200 35.900 ;
        RECT 181.400 32.100 181.800 37.900 ;
        RECT 182.200 34.700 182.600 35.100 ;
        RECT 182.200 29.200 182.500 34.700 ;
        RECT 171.000 26.100 171.400 26.200 ;
        RECT 171.800 26.100 172.200 26.200 ;
        RECT 171.000 25.800 172.200 26.100 ;
        RECT 174.200 25.900 174.600 26.300 ;
        RECT 175.000 23.100 175.400 28.900 ;
        RECT 177.400 28.800 177.800 29.200 ;
        RECT 178.200 29.100 178.600 29.200 ;
        RECT 179.000 29.100 179.400 29.200 ;
        RECT 178.200 28.800 179.400 29.100 ;
        RECT 177.400 28.200 177.700 28.800 ;
        RECT 176.600 25.100 177.000 27.900 ;
        RECT 177.400 27.800 177.800 28.200 ;
        RECT 177.400 19.200 177.700 27.800 ;
        RECT 179.000 25.800 179.400 26.200 ;
        RECT 173.400 19.100 173.800 19.200 ;
        RECT 174.200 19.100 174.600 19.200 ;
        RECT 173.400 18.800 174.600 19.100 ;
        RECT 177.400 18.800 177.800 19.200 ;
        RECT 168.600 15.800 169.000 16.200 ;
        RECT 175.800 16.100 176.200 16.200 ;
        RECT 176.600 16.100 177.000 16.200 ;
        RECT 175.800 15.800 177.000 16.100 ;
        RECT 178.200 15.800 178.600 16.200 ;
        RECT 168.600 15.200 168.900 15.800 ;
        RECT 168.600 14.800 169.000 15.200 ;
        RECT 171.000 14.800 171.400 15.200 ;
        RECT 172.600 15.100 173.000 15.200 ;
        RECT 173.400 15.100 173.800 15.200 ;
        RECT 172.600 14.800 173.800 15.100 ;
        RECT 169.400 13.800 169.800 14.200 ;
        RECT 170.200 13.800 170.600 14.200 ;
        RECT 167.000 12.100 167.400 12.200 ;
        RECT 167.800 12.100 168.200 12.200 ;
        RECT 167.000 11.800 168.200 12.100 ;
        RECT 168.600 11.800 169.000 12.200 ;
        RECT 167.000 8.800 167.400 9.200 ;
        RECT 161.400 5.100 161.800 7.900 ;
        RECT 162.200 7.800 162.600 8.200 ;
        RECT 163.000 7.800 163.400 8.200 ;
        RECT 167.000 7.200 167.300 8.800 ;
        RECT 167.000 6.800 167.400 7.200 ;
        RECT 163.000 6.100 163.400 6.200 ;
        RECT 163.800 6.100 164.200 6.200 ;
        RECT 163.000 5.800 164.200 6.100 ;
        RECT 167.000 6.100 167.400 6.200 ;
        RECT 167.800 6.100 168.200 6.200 ;
        RECT 168.600 6.100 168.900 11.800 ;
        RECT 167.000 5.800 168.900 6.100 ;
        RECT 169.400 5.200 169.700 13.800 ;
        RECT 170.200 12.200 170.500 13.800 ;
        RECT 170.200 11.800 170.600 12.200 ;
        RECT 171.000 6.100 171.300 14.800 ;
        RECT 178.200 14.200 178.500 15.800 ;
        RECT 179.000 15.200 179.300 25.800 ;
        RECT 179.800 25.100 180.200 27.900 ;
        RECT 180.600 26.800 181.000 27.200 ;
        RECT 180.600 26.200 180.900 26.800 ;
        RECT 180.600 25.800 181.000 26.200 ;
        RECT 181.400 23.100 181.800 28.900 ;
        RECT 182.200 28.800 182.600 29.200 ;
        RECT 182.200 26.300 182.500 28.800 ;
        RECT 182.200 25.900 182.600 26.300 ;
        RECT 182.200 25.800 182.500 25.900 ;
        RECT 183.000 25.100 183.300 53.800 ;
        RECT 183.800 53.100 184.200 55.900 ;
        RECT 185.400 52.100 185.800 57.900 ;
        RECT 186.200 56.800 186.600 57.200 ;
        RECT 186.200 55.100 186.500 56.800 ;
        RECT 186.200 54.700 186.600 55.100 ;
        RECT 187.000 54.200 187.300 63.800 ;
        RECT 192.600 59.200 192.900 69.800 ;
        RECT 193.400 69.200 193.700 71.800 ;
        RECT 193.400 68.800 193.800 69.200 ;
        RECT 193.400 59.800 193.800 60.200 ;
        RECT 193.400 59.200 193.700 59.800 ;
        RECT 192.600 58.800 193.000 59.200 ;
        RECT 193.400 58.800 193.800 59.200 ;
        RECT 187.000 53.800 187.400 54.200 ;
        RECT 190.200 52.100 190.600 57.900 ;
        RECT 191.000 52.800 191.400 53.200 ;
        RECT 193.400 53.100 193.800 53.200 ;
        RECT 194.200 53.100 194.600 53.200 ;
        RECT 193.400 52.800 194.600 53.100 ;
        RECT 191.000 49.200 191.300 52.800 ;
        RECT 183.800 43.100 184.200 48.900 ;
        RECT 185.400 46.800 185.800 47.200 ;
        RECT 185.400 46.200 185.700 46.800 ;
        RECT 184.600 45.800 185.000 46.200 ;
        RECT 185.400 45.800 185.800 46.200 ;
        RECT 187.000 45.800 187.400 46.200 ;
        RECT 182.200 24.800 183.300 25.100 ;
        RECT 179.800 15.800 180.200 16.200 ;
        RECT 179.800 15.200 180.100 15.800 ;
        RECT 179.000 14.800 179.400 15.200 ;
        RECT 179.800 14.800 180.200 15.200 ;
        RECT 181.400 14.800 181.800 15.200 ;
        RECT 177.400 13.800 177.800 14.200 ;
        RECT 178.200 13.800 178.600 14.200 ;
        RECT 180.600 13.800 181.000 14.200 ;
        RECT 177.400 12.200 177.700 13.800 ;
        RECT 180.600 12.200 180.900 13.800 ;
        RECT 181.400 13.200 181.700 14.800 ;
        RECT 181.400 12.800 181.800 13.200 ;
        RECT 172.600 11.800 173.000 12.200 ;
        RECT 175.800 11.800 176.200 12.200 ;
        RECT 177.400 11.800 177.800 12.200 ;
        RECT 180.600 11.800 181.000 12.200 ;
        RECT 172.600 9.200 172.900 11.800 ;
        RECT 175.800 9.200 176.100 11.800 ;
        RECT 172.600 8.800 173.000 9.200 ;
        RECT 171.800 7.800 172.200 8.200 ;
        RECT 171.800 7.200 172.100 7.800 ;
        RECT 171.800 6.800 172.200 7.200 ;
        RECT 171.800 6.100 172.200 6.200 ;
        RECT 171.000 5.800 172.200 6.100 ;
        RECT 163.000 4.800 163.400 5.200 ;
        RECT 169.400 4.800 169.800 5.200 ;
        RECT 163.000 4.200 163.300 4.800 ;
        RECT 163.000 3.800 163.400 4.200 ;
        RECT 175.000 3.100 175.400 8.900 ;
        RECT 175.800 8.800 176.200 9.200 ;
        RECT 178.200 7.800 178.600 8.200 ;
        RECT 175.800 6.800 176.200 7.200 ;
        RECT 175.800 6.200 176.100 6.800 ;
        RECT 178.200 6.200 178.500 7.800 ;
        RECT 175.800 5.800 176.200 6.200 ;
        RECT 178.200 5.800 178.600 6.200 ;
        RECT 179.800 3.100 180.200 8.900 ;
        RECT 182.200 8.200 182.500 24.800 ;
        RECT 184.600 19.200 184.900 45.800 ;
        RECT 186.200 32.100 186.600 37.900 ;
        RECT 187.000 37.200 187.300 45.800 ;
        RECT 188.600 43.100 189.000 48.900 ;
        RECT 191.000 48.800 191.400 49.200 ;
        RECT 187.000 36.800 187.400 37.200 ;
        RECT 186.200 23.100 186.600 28.900 ;
        RECT 184.600 18.800 185.000 19.200 ;
        RECT 187.000 19.100 187.300 36.800 ;
        RECT 188.600 31.800 189.000 32.200 ;
        RECT 188.600 29.200 188.900 31.800 ;
        RECT 188.600 28.800 189.000 29.200 ;
        RECT 186.200 18.800 187.300 19.100 ;
        RECT 188.600 21.800 189.000 22.200 ;
        RECT 183.000 15.100 183.400 15.200 ;
        RECT 183.800 15.100 184.200 15.200 ;
        RECT 183.000 14.800 184.200 15.100 ;
        RECT 183.800 13.800 184.200 14.200 ;
        RECT 183.800 13.200 184.100 13.800 ;
        RECT 183.000 12.800 183.400 13.200 ;
        RECT 183.800 12.800 184.200 13.200 ;
        RECT 185.400 13.100 185.800 15.900 ;
        RECT 186.200 14.200 186.500 18.800 ;
        RECT 186.200 13.800 186.600 14.200 ;
        RECT 183.000 12.200 183.300 12.800 ;
        RECT 183.000 11.800 183.400 12.200 ;
        RECT 183.800 8.200 184.100 12.800 ;
        RECT 187.000 12.100 187.400 17.900 ;
        RECT 188.600 16.200 188.900 21.800 ;
        RECT 188.600 15.800 189.000 16.200 ;
        RECT 187.800 14.700 188.200 15.200 ;
        RECT 181.400 5.100 181.800 7.900 ;
        RECT 182.200 7.800 182.600 8.200 ;
        RECT 183.800 7.800 184.200 8.200 ;
        RECT 182.200 5.800 182.600 6.200 ;
        RECT 182.200 5.200 182.500 5.800 ;
        RECT 182.200 4.800 182.600 5.200 ;
        RECT 184.600 5.100 185.000 7.900 ;
        RECT 185.400 7.800 185.800 8.200 ;
        RECT 185.400 7.200 185.700 7.800 ;
        RECT 185.400 6.800 185.800 7.200 ;
        RECT 186.200 3.100 186.600 8.900 ;
        RECT 187.800 6.200 188.100 14.700 ;
        RECT 191.800 12.100 192.200 17.900 ;
        RECT 194.200 12.800 194.600 13.200 ;
        RECT 194.200 12.200 194.500 12.800 ;
        RECT 194.200 11.800 194.600 12.200 ;
        RECT 194.200 9.200 194.500 11.800 ;
        RECT 187.800 5.800 188.200 6.200 ;
        RECT 191.000 3.100 191.400 8.900 ;
        RECT 194.200 8.800 194.600 9.200 ;
      LAYER via2 ;
        RECT 20.600 167.800 21.000 168.200 ;
        RECT 8.600 165.800 9.000 166.200 ;
        RECT 16.600 165.800 17.000 166.200 ;
        RECT 1.400 143.800 1.800 144.200 ;
        RECT 1.400 123.800 1.800 124.200 ;
        RECT 23.800 161.800 24.200 162.200 ;
        RECT 43.000 167.800 43.400 168.200 ;
        RECT 18.200 141.800 18.600 142.200 ;
        RECT 30.200 151.800 30.600 152.200 ;
        RECT 12.600 114.800 13.000 115.200 ;
        RECT 14.200 114.000 14.600 114.400 ;
        RECT 7.800 107.800 8.200 108.200 ;
        RECT 1.400 106.800 1.800 107.200 ;
        RECT 1.400 86.800 1.800 87.200 ;
        RECT 14.200 98.800 14.600 99.200 ;
        RECT 7.800 92.800 8.200 93.200 ;
        RECT 3.800 48.800 4.200 49.200 ;
        RECT 1.400 38.800 1.800 39.200 ;
        RECT 24.600 132.800 25.000 133.200 ;
        RECT 30.200 134.800 30.600 135.200 ;
        RECT 41.400 154.800 41.800 155.200 ;
        RECT 51.800 161.800 52.200 162.200 ;
        RECT 52.600 151.800 53.000 152.200 ;
        RECT 37.400 144.800 37.800 145.200 ;
        RECT 33.400 125.800 33.800 126.200 ;
        RECT 51.800 146.800 52.200 147.200 ;
        RECT 63.000 147.800 63.400 148.200 ;
        RECT 55.800 144.800 56.200 145.200 ;
        RECT 42.200 133.800 42.600 134.200 ;
        RECT 35.800 113.800 36.200 114.200 ;
        RECT 23.800 106.800 24.200 107.200 ;
        RECT 19.800 104.800 20.200 105.200 ;
        RECT 35.000 105.800 35.400 106.200 ;
        RECT 16.600 74.800 17.000 75.200 ;
        RECT 26.200 93.800 26.600 94.200 ;
        RECT 30.200 92.800 30.600 93.200 ;
        RECT 51.800 116.800 52.200 117.200 ;
        RECT 55.800 125.800 56.200 126.200 ;
        RECT 71.800 144.800 72.200 145.200 ;
        RECT 75.000 141.800 75.400 142.200 ;
        RECT 87.000 165.800 87.400 166.200 ;
        RECT 89.400 165.800 89.800 166.200 ;
        RECT 87.000 154.800 87.400 155.200 ;
        RECT 79.800 145.900 80.200 146.300 ;
        RECT 66.200 136.800 66.600 137.200 ;
        RECT 59.800 127.800 60.200 128.200 ;
        RECT 37.400 107.800 37.800 108.200 ;
        RECT 54.200 114.800 54.600 115.200 ;
        RECT 67.800 134.800 68.200 135.200 ;
        RECT 74.200 136.800 74.600 137.200 ;
        RECT 59.000 123.800 59.400 124.200 ;
        RECT 59.800 115.800 60.200 116.200 ;
        RECT 42.200 103.800 42.600 104.200 ;
        RECT 33.400 93.800 33.800 94.200 ;
        RECT 47.800 105.800 48.200 106.200 ;
        RECT 47.000 94.800 47.400 95.200 ;
        RECT 32.600 87.800 33.000 88.200 ;
        RECT 28.600 86.800 29.000 87.200 ;
        RECT 35.800 84.800 36.200 85.200 ;
        RECT 44.600 86.800 45.000 87.200 ;
        RECT 84.600 147.800 85.000 148.200 ;
        RECT 91.800 161.800 92.200 162.200 ;
        RECT 107.800 161.800 108.200 162.200 ;
        RECT 99.000 156.800 99.400 157.200 ;
        RECT 102.200 154.800 102.600 155.200 ;
        RECT 108.600 154.800 109.000 155.200 ;
        RECT 126.200 154.800 126.600 155.200 ;
        RECT 104.600 148.800 105.000 149.200 ;
        RECT 87.000 145.800 87.400 146.200 ;
        RECT 78.200 123.800 78.600 124.200 ;
        RECT 59.800 104.800 60.200 105.200 ;
        RECT 59.800 94.800 60.200 95.200 ;
        RECT 83.000 128.800 83.400 129.200 ;
        RECT 83.000 124.800 83.400 125.200 ;
        RECT 85.400 125.800 85.800 126.200 ;
        RECT 86.200 113.800 86.600 114.200 ;
        RECT 93.400 134.800 93.800 135.200 ;
        RECT 91.800 133.800 92.200 134.200 ;
        RECT 93.400 112.800 93.800 113.200 ;
        RECT 64.600 105.800 65.000 106.200 ;
        RECT 66.200 105.800 66.600 106.200 ;
        RECT 67.800 105.800 68.200 106.200 ;
        RECT 59.000 92.800 59.400 93.200 ;
        RECT 63.000 88.800 63.400 89.200 ;
        RECT 60.600 85.800 61.000 86.200 ;
        RECT 47.800 72.800 48.200 73.200 ;
        RECT 50.200 72.800 50.600 73.200 ;
        RECT 51.800 72.800 52.200 73.200 ;
        RECT 43.000 48.800 43.400 49.200 ;
        RECT 24.600 33.800 25.000 34.200 ;
        RECT 7.800 23.800 8.200 24.200 ;
        RECT 3.800 11.800 4.200 12.200 ;
        RECT 12.600 25.800 13.000 26.200 ;
        RECT 30.200 31.800 30.600 32.200 ;
        RECT 48.600 48.800 49.000 49.200 ;
        RECT 18.200 21.800 18.600 22.200 ;
        RECT 12.600 8.800 13.000 9.200 ;
        RECT 13.400 7.800 13.800 8.200 ;
        RECT 40.600 34.800 41.000 35.200 ;
        RECT 45.400 34.800 45.800 35.200 ;
        RECT 38.200 25.800 38.600 26.200 ;
        RECT 53.400 32.800 53.800 33.200 ;
        RECT 80.600 92.800 81.000 93.200 ;
        RECT 87.800 92.800 88.200 93.200 ;
        RECT 122.200 153.800 122.600 154.200 ;
        RECT 123.800 147.800 124.200 148.200 ;
        RECT 151.000 165.800 151.400 166.200 ;
        RECT 155.000 161.800 155.400 162.200 ;
        RECT 151.800 152.800 152.200 153.200 ;
        RECT 161.400 146.800 161.800 147.200 ;
        RECT 163.000 144.800 163.400 145.200 ;
        RECT 166.200 144.800 166.600 145.200 ;
        RECT 105.400 134.800 105.800 135.200 ;
        RECT 123.800 134.800 124.200 135.200 ;
        RECT 81.400 75.800 81.800 76.200 ;
        RECT 81.400 74.800 81.800 75.200 ;
        RECT 80.600 73.800 81.000 74.200 ;
        RECT 79.800 72.800 80.200 73.200 ;
        RECT 136.600 134.800 137.000 135.200 ;
        RECT 138.200 134.800 138.600 135.200 ;
        RECT 145.400 131.800 145.800 132.200 ;
        RECT 160.600 132.800 161.000 133.200 ;
        RECT 85.400 74.800 85.800 75.200 ;
        RECT 86.200 73.800 86.600 74.200 ;
        RECT 119.800 97.800 120.200 98.200 ;
        RECT 117.400 93.800 117.800 94.200 ;
        RECT 87.800 67.800 88.200 68.200 ;
        RECT 87.800 65.800 88.200 66.200 ;
        RECT 94.200 66.800 94.600 67.200 ;
        RECT 146.200 125.800 146.600 126.200 ;
        RECT 131.000 114.800 131.400 115.200 ;
        RECT 131.000 93.800 131.400 94.200 ;
        RECT 126.200 85.800 126.600 86.200 ;
        RECT 126.200 74.800 126.600 75.200 ;
        RECT 127.800 72.800 128.200 73.200 ;
        RECT 159.000 124.800 159.400 125.200 ;
        RECT 156.600 105.800 157.000 106.200 ;
        RECT 139.800 91.800 140.200 92.200 ;
        RECT 162.200 125.800 162.600 126.200 ;
        RECT 167.800 133.800 168.200 134.200 ;
        RECT 172.600 134.800 173.000 135.200 ;
        RECT 163.000 107.800 163.400 108.200 ;
        RECT 162.200 106.800 162.600 107.200 ;
        RECT 167.800 106.800 168.200 107.200 ;
        RECT 184.600 134.800 185.000 135.200 ;
        RECT 191.800 125.800 192.200 126.200 ;
        RECT 185.400 114.800 185.800 115.200 ;
        RECT 186.200 94.700 186.600 95.100 ;
        RECT 163.800 86.800 164.200 87.200 ;
        RECT 165.400 85.800 165.800 86.200 ;
        RECT 135.000 65.800 135.400 66.200 ;
        RECT 159.000 74.800 159.400 75.200 ;
        RECT 168.600 83.800 169.000 84.200 ;
        RECT 171.000 83.800 171.400 84.200 ;
        RECT 168.600 75.800 169.000 76.200 ;
        RECT 169.400 72.800 169.800 73.200 ;
        RECT 167.800 71.800 168.200 72.200 ;
        RECT 155.000 66.800 155.400 67.200 ;
        RECT 163.000 66.800 163.400 67.200 ;
        RECT 154.200 65.800 154.600 66.200 ;
        RECT 83.800 55.800 84.200 56.200 ;
        RECT 108.600 54.800 109.000 55.200 ;
        RECT 68.600 47.800 69.000 48.200 ;
        RECT 79.000 48.800 79.400 49.200 ;
        RECT 82.200 46.800 82.600 47.200 ;
        RECT 72.600 33.800 73.000 34.200 ;
        RECT 23.000 6.800 23.400 7.200 ;
        RECT 3.800 5.800 4.200 6.200 ;
        RECT 5.400 4.800 5.800 5.200 ;
        RECT 19.800 4.800 20.200 5.200 ;
        RECT 35.800 8.800 36.200 9.200 ;
        RECT 59.800 13.800 60.200 14.200 ;
        RECT 79.000 32.800 79.400 33.200 ;
        RECT 75.000 25.800 75.400 26.200 ;
        RECT 77.400 25.800 77.800 26.200 ;
        RECT 91.000 44.800 91.400 45.200 ;
        RECT 88.600 38.800 89.000 39.200 ;
        RECT 85.400 34.800 85.800 35.200 ;
        RECT 75.800 23.800 76.200 24.200 ;
        RECT 98.200 51.800 98.600 52.200 ;
        RECT 100.600 48.800 101.000 49.200 ;
        RECT 79.000 21.800 79.400 22.200 ;
        RECT 55.000 4.800 55.400 5.200 ;
        RECT 114.200 54.800 114.600 55.200 ;
        RECT 103.800 33.800 104.200 34.200 ;
        RECT 81.400 13.800 81.800 14.200 ;
        RECT 91.800 13.800 92.200 14.200 ;
        RECT 77.400 6.800 77.800 7.200 ;
        RECT 87.800 4.800 88.200 5.200 ;
        RECT 107.800 13.800 108.200 14.200 ;
        RECT 103.800 8.800 104.200 9.200 ;
        RECT 133.400 45.800 133.800 46.200 ;
        RECT 139.800 48.800 140.200 49.200 ;
        RECT 145.400 54.800 145.800 55.200 ;
        RECT 153.400 47.800 153.800 48.200 ;
        RECT 159.000 48.800 159.400 49.200 ;
        RECT 155.000 45.800 155.400 46.200 ;
        RECT 157.400 45.800 157.800 46.200 ;
        RECT 156.600 43.800 157.000 44.200 ;
        RECT 151.800 34.800 152.200 35.200 ;
        RECT 123.000 7.800 123.400 8.200 ;
        RECT 134.200 15.800 134.600 16.200 ;
        RECT 139.800 15.800 140.200 16.200 ;
        RECT 127.000 5.800 127.400 6.200 ;
        RECT 126.200 4.800 126.600 5.200 ;
        RECT 149.400 25.800 149.800 26.200 ;
        RECT 155.000 28.800 155.400 29.200 ;
        RECT 174.200 65.800 174.600 66.200 ;
        RECT 175.800 54.800 176.200 55.200 ;
        RECT 177.400 54.800 177.800 55.200 ;
        RECT 179.000 53.800 179.400 54.200 ;
        RECT 169.400 47.800 169.800 48.200 ;
        RECT 171.000 45.800 171.400 46.200 ;
        RECT 168.600 44.800 169.000 45.200 ;
        RECT 168.600 34.800 169.000 35.200 ;
        RECT 155.000 13.800 155.400 14.200 ;
        RECT 165.400 28.800 165.800 29.200 ;
        RECT 171.800 25.800 172.200 26.200 ;
        RECT 179.000 28.800 179.400 29.200 ;
        RECT 176.600 15.800 177.000 16.200 ;
        RECT 167.800 5.800 168.200 6.200 ;
        RECT 183.800 14.800 184.200 15.200 ;
        RECT 187.800 14.800 188.200 15.200 ;
      LAYER metal3 ;
        RECT 6.200 167.800 6.600 168.200 ;
        RECT 9.400 168.100 9.800 168.200 ;
        RECT 12.600 168.100 13.000 168.200 ;
        RECT 9.400 167.800 13.000 168.100 ;
        RECT 13.400 167.800 13.800 168.200 ;
        RECT 20.600 168.100 21.000 168.200 ;
        RECT 21.400 168.100 21.800 168.200 ;
        RECT 20.600 167.800 21.800 168.100 ;
        RECT 40.600 168.100 41.000 168.200 ;
        RECT 43.000 168.100 43.400 168.200 ;
        RECT 62.200 168.100 62.600 168.200 ;
        RECT 40.600 167.800 62.600 168.100 ;
        RECT 115.000 168.100 115.400 168.200 ;
        RECT 138.200 168.100 138.600 168.200 ;
        RECT 144.600 168.100 145.000 168.200 ;
        RECT 115.000 167.800 145.000 168.100 ;
        RECT 2.200 167.100 2.600 167.200 ;
        RECT 6.200 167.100 6.500 167.800 ;
        RECT 2.200 166.800 6.500 167.100 ;
        RECT 11.000 167.100 11.400 167.200 ;
        RECT 13.400 167.100 13.700 167.800 ;
        RECT 18.200 167.100 18.600 167.200 ;
        RECT 11.000 166.800 12.900 167.100 ;
        RECT 13.400 166.800 18.600 167.100 ;
        RECT 43.000 166.800 43.400 167.200 ;
        RECT 43.800 166.800 44.200 167.200 ;
        RECT 57.400 166.800 57.800 167.200 ;
        RECT 62.200 167.100 62.600 167.200 ;
        RECT 69.400 167.100 69.800 167.200 ;
        RECT 62.200 166.800 69.800 167.100 ;
        RECT 97.400 166.800 97.800 167.200 ;
        RECT 127.000 167.100 127.400 167.200 ;
        RECT 139.000 167.100 139.400 167.200 ;
        RECT 145.400 167.100 145.800 167.200 ;
        RECT 127.000 166.800 145.800 167.100 ;
        RECT 147.000 167.100 147.400 167.200 ;
        RECT 151.000 167.100 151.400 167.200 ;
        RECT 147.000 166.800 151.400 167.100 ;
        RECT 159.800 166.800 160.200 167.200 ;
        RECT 5.400 166.100 5.800 166.200 ;
        RECT 8.600 166.100 9.000 166.200 ;
        RECT 5.400 165.800 9.000 166.100 ;
        RECT 11.800 165.800 12.200 166.200 ;
        RECT 12.600 166.100 12.900 166.800 ;
        RECT 16.600 166.100 17.000 166.200 ;
        RECT 43.000 166.100 43.300 166.800 ;
        RECT 12.600 165.800 17.000 166.100 ;
        RECT 29.400 165.800 43.300 166.100 ;
        RECT 43.800 166.100 44.100 166.800 ;
        RECT 47.800 166.100 48.200 166.200 ;
        RECT 57.400 166.100 57.700 166.800 ;
        RECT 61.400 166.100 61.800 166.200 ;
        RECT 66.200 166.100 66.600 166.200 ;
        RECT 43.800 165.800 48.900 166.100 ;
        RECT 57.400 165.800 66.600 166.100 ;
        RECT 87.000 166.100 87.400 166.200 ;
        RECT 89.400 166.100 89.800 166.200 ;
        RECT 87.000 165.800 89.800 166.100 ;
        RECT 97.400 166.100 97.700 166.800 ;
        RECT 100.600 166.100 101.000 166.200 ;
        RECT 111.800 166.100 112.200 166.200 ;
        RECT 97.400 165.800 112.200 166.100 ;
        RECT 144.600 166.100 145.000 166.200 ;
        RECT 151.000 166.100 151.400 166.200 ;
        RECT 144.600 165.800 151.400 166.100 ;
        RECT 159.800 166.100 160.100 166.800 ;
        RECT 167.000 166.100 167.400 166.200 ;
        RECT 179.000 166.100 179.400 166.200 ;
        RECT 159.800 165.800 167.400 166.100 ;
        RECT 169.400 165.800 179.400 166.100 ;
        RECT 11.800 165.100 12.100 165.800 ;
        RECT 29.400 165.200 29.700 165.800 ;
        RECT 39.000 165.200 39.300 165.800 ;
        RECT 169.400 165.200 169.700 165.800 ;
        RECT 15.000 165.100 15.400 165.200 ;
        RECT 11.800 164.800 15.400 165.100 ;
        RECT 29.400 164.800 29.800 165.200 ;
        RECT 39.000 164.800 39.400 165.200 ;
        RECT 49.400 165.100 49.800 165.200 ;
        RECT 72.600 165.100 73.000 165.200 ;
        RECT 49.400 164.800 73.000 165.100 ;
        RECT 102.200 164.800 102.600 165.200 ;
        RECT 103.800 165.100 104.200 165.200 ;
        RECT 111.800 165.100 112.200 165.200 ;
        RECT 103.800 164.800 112.200 165.100 ;
        RECT 169.400 164.800 169.800 165.200 ;
        RECT 102.200 164.200 102.500 164.800 ;
        RECT 7.000 164.100 7.400 164.200 ;
        RECT 10.200 164.100 10.600 164.200 ;
        RECT 14.200 164.100 14.600 164.200 ;
        RECT 26.200 164.100 26.600 164.200 ;
        RECT 7.000 163.800 26.600 164.100 ;
        RECT 60.600 164.100 61.000 164.200 ;
        RECT 64.600 164.100 65.000 164.200 ;
        RECT 60.600 163.800 65.000 164.100 ;
        RECT 102.200 163.800 102.600 164.200 ;
        RECT 163.000 164.100 163.400 164.200 ;
        RECT 192.600 164.100 193.000 164.200 ;
        RECT 163.000 163.800 193.000 164.100 ;
        RECT 80.600 163.100 81.000 163.200 ;
        RECT 82.200 163.100 82.600 163.200 ;
        RECT 94.200 163.100 94.600 163.200 ;
        RECT 80.600 162.800 94.600 163.100 ;
        RECT 124.600 162.800 125.000 163.200 ;
        RECT 124.600 162.200 124.900 162.800 ;
        RECT 23.800 162.100 24.200 162.200 ;
        RECT 25.400 162.100 25.800 162.200 ;
        RECT 31.800 162.100 32.200 162.200 ;
        RECT 47.000 162.100 47.400 162.200 ;
        RECT 23.800 161.800 47.400 162.100 ;
        RECT 51.800 162.100 52.200 162.200 ;
        RECT 63.000 162.100 63.400 162.200 ;
        RECT 51.800 161.800 63.400 162.100 ;
        RECT 86.200 162.100 86.600 162.200 ;
        RECT 91.800 162.100 92.200 162.200 ;
        RECT 107.800 162.100 108.200 162.200 ;
        RECT 111.000 162.100 111.400 162.200 ;
        RECT 86.200 161.800 111.400 162.100 ;
        RECT 124.600 161.800 125.000 162.200 ;
        RECT 155.000 162.100 155.400 162.200 ;
        RECT 165.400 162.100 165.800 162.200 ;
        RECT 155.000 161.800 165.800 162.100 ;
        RECT 119.000 160.100 119.400 160.200 ;
        RECT 127.000 160.100 127.400 160.200 ;
        RECT 129.400 160.100 129.800 160.200 ;
        RECT 119.000 159.800 129.800 160.100 ;
        RECT 56.600 159.100 57.000 159.200 ;
        RECT 147.800 159.100 148.200 159.200 ;
        RECT 161.400 159.100 161.800 159.200 ;
        RECT 56.600 158.800 161.800 159.100 ;
        RECT 43.800 158.100 44.200 158.200 ;
        RECT 44.600 158.100 45.000 158.200 ;
        RECT 43.800 157.800 45.000 158.100 ;
        RECT 121.400 158.100 121.800 158.200 ;
        RECT 131.000 158.100 131.400 158.200 ;
        RECT 144.600 158.100 145.000 158.200 ;
        RECT 121.400 157.800 145.000 158.100 ;
        RECT 175.800 158.100 176.200 158.200 ;
        RECT 191.000 158.100 191.400 158.200 ;
        RECT 175.800 157.800 191.400 158.100 ;
        RECT 99.000 157.100 99.400 157.200 ;
        RECT 103.000 157.100 103.400 157.200 ;
        RECT 99.000 156.800 103.400 157.100 ;
        RECT 35.800 155.800 36.200 156.200 ;
        RECT 37.400 156.100 37.800 156.200 ;
        RECT 55.000 156.100 55.400 156.200 ;
        RECT 37.400 155.800 55.400 156.100 ;
        RECT 72.600 156.100 73.000 156.200 ;
        RECT 91.000 156.100 91.400 156.200 ;
        RECT 72.600 155.800 91.400 156.100 ;
        RECT 95.000 156.100 95.400 156.200 ;
        RECT 101.400 156.100 101.800 156.200 ;
        RECT 95.000 155.800 101.800 156.100 ;
        RECT 118.200 156.100 118.600 156.200 ;
        RECT 123.800 156.100 124.200 156.200 ;
        RECT 118.200 155.800 124.200 156.100 ;
        RECT 128.600 155.800 129.000 156.200 ;
        RECT 146.200 155.800 146.600 156.200 ;
        RECT 151.000 155.800 151.400 156.200 ;
        RECT 185.400 155.800 185.800 156.200 ;
        RECT 16.600 155.100 17.000 155.200 ;
        RECT 19.800 155.100 20.200 155.200 ;
        RECT 16.600 154.800 20.200 155.100 ;
        RECT 35.800 155.100 36.100 155.800 ;
        RECT 41.400 155.100 41.800 155.200 ;
        RECT 87.000 155.100 87.400 155.200 ;
        RECT 35.800 154.800 41.800 155.100 ;
        RECT 77.400 154.800 87.400 155.100 ;
        RECT 95.800 155.100 96.200 155.200 ;
        RECT 99.800 155.100 100.200 155.200 ;
        RECT 95.800 154.800 100.200 155.100 ;
        RECT 102.200 155.100 102.600 155.200 ;
        RECT 108.600 155.100 109.000 155.200 ;
        RECT 102.200 154.800 109.000 155.100 ;
        RECT 115.000 155.100 115.400 155.200 ;
        RECT 121.400 155.100 121.800 155.200 ;
        RECT 115.000 154.800 121.800 155.100 ;
        RECT 126.200 155.100 126.600 155.200 ;
        RECT 127.800 155.100 128.200 155.200 ;
        RECT 126.200 154.800 128.200 155.100 ;
        RECT 128.600 155.100 128.900 155.800 ;
        RECT 134.200 155.100 134.600 155.200 ;
        RECT 139.000 155.100 139.400 155.200 ;
        RECT 139.800 155.100 140.200 155.200 ;
        RECT 128.600 154.800 130.500 155.100 ;
        RECT 134.200 154.800 140.200 155.100 ;
        RECT 146.200 155.100 146.500 155.800 ;
        RECT 151.000 155.100 151.300 155.800 ;
        RECT 146.200 154.800 151.300 155.100 ;
        RECT 154.200 154.800 154.600 155.200 ;
        RECT 174.200 155.100 174.600 155.200 ;
        RECT 175.800 155.100 176.200 155.200 ;
        RECT 174.200 154.800 176.200 155.100 ;
        RECT 181.400 155.100 181.800 155.200 ;
        RECT 185.400 155.100 185.700 155.800 ;
        RECT 181.400 154.800 185.700 155.100 ;
        RECT 77.400 154.200 77.700 154.800 ;
        RECT 14.200 154.100 14.600 154.200 ;
        RECT 19.000 154.100 19.400 154.200 ;
        RECT 23.800 154.100 24.200 154.200 ;
        RECT 28.600 154.100 29.000 154.200 ;
        RECT 51.000 154.100 51.400 154.200 ;
        RECT 60.600 154.100 61.000 154.200 ;
        RECT 14.200 153.800 51.400 154.100 ;
        RECT 59.800 153.800 61.000 154.100 ;
        RECT 77.400 153.800 77.800 154.200 ;
        RECT 84.600 154.100 85.000 154.200 ;
        RECT 92.600 154.100 93.000 154.200 ;
        RECT 95.800 154.100 96.100 154.800 ;
        RECT 84.600 153.800 96.100 154.100 ;
        RECT 122.200 154.100 122.600 154.200 ;
        RECT 126.200 154.100 126.500 154.800 ;
        RECT 122.200 153.800 126.500 154.100 ;
        RECT 130.200 154.200 130.500 154.800 ;
        RECT 130.200 153.800 130.600 154.200 ;
        RECT 144.600 154.100 145.000 154.200 ;
        RECT 152.600 154.100 153.000 154.200 ;
        RECT 154.200 154.100 154.500 154.800 ;
        RECT 174.200 154.200 174.500 154.800 ;
        RECT 166.200 154.100 166.600 154.200 ;
        RECT 144.600 153.800 166.600 154.100 ;
        RECT 174.200 153.800 174.600 154.200 ;
        RECT 177.400 154.100 177.800 154.200 ;
        RECT 180.600 154.100 181.000 154.200 ;
        RECT 177.400 153.800 181.000 154.100 ;
        RECT 59.800 153.200 60.100 153.800 ;
        RECT 59.800 152.800 60.200 153.200 ;
        RECT 69.400 153.100 69.800 153.200 ;
        RECT 77.400 153.100 77.800 153.200 ;
        RECT 69.400 152.800 77.800 153.100 ;
        RECT 90.200 153.100 90.600 153.200 ;
        RECT 95.800 153.100 96.200 153.200 ;
        RECT 96.600 153.100 97.000 153.200 ;
        RECT 90.200 152.800 97.000 153.100 ;
        RECT 101.400 153.100 101.800 153.200 ;
        RECT 103.800 153.100 104.200 153.200 ;
        RECT 101.400 152.800 104.200 153.100 ;
        RECT 108.600 153.100 109.000 153.200 ;
        RECT 119.000 153.100 119.400 153.200 ;
        RECT 108.600 152.800 119.400 153.100 ;
        RECT 129.400 153.100 129.800 153.200 ;
        RECT 132.600 153.100 133.000 153.200 ;
        RECT 129.400 152.800 133.000 153.100 ;
        RECT 134.200 153.100 134.600 153.200 ;
        RECT 138.200 153.100 138.600 153.200 ;
        RECT 134.200 152.800 138.600 153.100 ;
        RECT 151.800 153.100 152.200 153.200 ;
        RECT 154.200 153.100 154.600 153.200 ;
        RECT 156.600 153.100 157.000 153.200 ;
        RECT 151.800 152.800 157.000 153.100 ;
        RECT 165.400 153.100 165.800 153.200 ;
        RECT 171.800 153.100 172.200 153.200 ;
        RECT 165.400 152.800 172.200 153.100 ;
        RECT 30.200 152.100 30.600 152.200 ;
        RECT 43.000 152.100 43.400 152.200 ;
        RECT 47.000 152.100 47.400 152.200 ;
        RECT 30.200 151.800 47.400 152.100 ;
        RECT 52.600 152.100 53.000 152.200 ;
        RECT 58.200 152.100 58.600 152.200 ;
        RECT 60.600 152.100 61.000 152.200 ;
        RECT 52.600 151.800 61.000 152.100 ;
        RECT 119.800 152.100 120.200 152.200 ;
        RECT 125.400 152.100 125.800 152.200 ;
        RECT 119.800 151.800 125.800 152.100 ;
        RECT 132.600 152.100 133.000 152.200 ;
        RECT 132.600 151.800 135.300 152.100 ;
        RECT 135.000 151.200 135.300 151.800 ;
        RECT 20.600 151.100 21.000 151.200 ;
        RECT 56.600 151.100 57.000 151.200 ;
        RECT 20.600 150.800 57.000 151.100 ;
        RECT 57.400 151.100 57.800 151.200 ;
        RECT 61.400 151.100 61.800 151.200 ;
        RECT 67.000 151.100 67.400 151.200 ;
        RECT 57.400 150.800 67.400 151.100 ;
        RECT 71.000 151.100 71.400 151.200 ;
        RECT 80.600 151.100 81.000 151.200 ;
        RECT 81.400 151.100 81.800 151.200 ;
        RECT 71.000 150.800 81.800 151.100 ;
        RECT 110.200 151.100 110.600 151.200 ;
        RECT 127.000 151.100 127.400 151.200 ;
        RECT 110.200 150.800 127.400 151.100 ;
        RECT 135.000 150.800 135.400 151.200 ;
        RECT 31.000 150.100 31.400 150.200 ;
        RECT 42.200 150.100 42.600 150.200 ;
        RECT 31.000 149.800 42.600 150.100 ;
        RECT 51.000 150.100 51.400 150.200 ;
        RECT 68.600 150.100 69.000 150.200 ;
        RECT 51.000 149.800 69.000 150.100 ;
        RECT 53.400 148.800 53.800 149.200 ;
        RECT 71.000 148.800 71.400 149.200 ;
        RECT 91.000 149.100 91.400 149.200 ;
        RECT 104.600 149.100 105.000 149.200 ;
        RECT 113.400 149.100 113.800 149.200 ;
        RECT 145.400 149.100 145.800 149.200 ;
        RECT 91.000 148.800 145.800 149.100 ;
        RECT 147.000 149.100 147.400 149.200 ;
        RECT 171.800 149.100 172.200 149.200 ;
        RECT 175.000 149.100 175.400 149.200 ;
        RECT 182.200 149.100 182.600 149.200 ;
        RECT 147.000 148.800 182.600 149.100 ;
        RECT 23.800 148.100 24.200 148.200 ;
        RECT 33.400 148.100 33.800 148.200 ;
        RECT 53.400 148.100 53.700 148.800 ;
        RECT 23.800 147.800 53.700 148.100 ;
        RECT 63.000 148.100 63.400 148.200 ;
        RECT 71.000 148.100 71.300 148.800 ;
        RECT 63.000 147.800 71.300 148.100 ;
        RECT 82.200 148.100 82.600 148.200 ;
        RECT 84.600 148.100 85.000 148.200 ;
        RECT 102.200 148.100 102.600 148.200 ;
        RECT 103.000 148.100 103.400 148.200 ;
        RECT 82.200 147.800 103.400 148.100 ;
        RECT 103.800 148.100 104.200 148.200 ;
        RECT 117.400 148.100 117.800 148.200 ;
        RECT 103.800 147.800 117.800 148.100 ;
        RECT 121.400 147.800 121.800 148.200 ;
        RECT 123.000 148.100 123.400 148.200 ;
        RECT 123.800 148.100 124.200 148.200 ;
        RECT 123.000 147.800 124.200 148.100 ;
        RECT 126.200 148.100 126.600 148.200 ;
        RECT 148.600 148.100 149.000 148.200 ;
        RECT 126.200 147.800 149.000 148.100 ;
        RECT 162.200 148.100 162.600 148.200 ;
        RECT 163.000 148.100 163.400 148.200 ;
        RECT 162.200 147.800 163.400 148.100 ;
        RECT 167.000 147.800 167.400 148.200 ;
        RECT 6.200 146.800 6.600 147.200 ;
        RECT 11.000 146.800 11.400 147.200 ;
        RECT 11.800 146.800 12.200 147.200 ;
        RECT 36.600 147.100 37.000 147.200 ;
        RECT 39.800 147.100 40.200 147.200 ;
        RECT 36.600 146.800 40.200 147.100 ;
        RECT 40.600 147.100 41.000 147.200 ;
        RECT 42.200 147.100 42.600 147.200 ;
        RECT 40.600 146.800 42.600 147.100 ;
        RECT 43.800 147.100 44.200 147.200 ;
        RECT 51.800 147.100 52.200 147.200 ;
        RECT 67.000 147.100 67.400 147.200 ;
        RECT 43.800 146.800 67.400 147.100 ;
        RECT 78.200 147.100 78.600 147.200 ;
        RECT 86.200 147.100 86.600 147.200 ;
        RECT 78.200 146.800 86.600 147.100 ;
        RECT 88.600 147.100 89.000 147.200 ;
        RECT 88.600 146.800 99.300 147.100 ;
        RECT 6.200 146.100 6.500 146.800 ;
        RECT 11.000 146.100 11.300 146.800 ;
        RECT 6.200 145.800 11.300 146.100 ;
        RECT 11.800 146.100 12.100 146.800 ;
        RECT 14.200 146.100 14.600 146.200 ;
        RECT 25.400 146.100 25.800 146.200 ;
        RECT 37.400 146.100 37.800 146.200 ;
        RECT 11.800 145.800 15.300 146.100 ;
        RECT 25.400 145.800 37.800 146.100 ;
        RECT 41.400 146.100 41.800 146.200 ;
        RECT 44.600 146.100 45.000 146.200 ;
        RECT 41.400 145.800 45.000 146.100 ;
        RECT 51.000 146.100 51.400 146.200 ;
        RECT 52.600 146.100 53.000 146.200 ;
        RECT 51.000 145.800 53.000 146.100 ;
        RECT 57.400 146.100 57.800 146.200 ;
        RECT 59.000 146.100 59.400 146.200 ;
        RECT 57.400 145.800 59.400 146.100 ;
        RECT 79.800 146.100 80.200 146.300 ;
        RECT 99.000 146.200 99.300 146.800 ;
        RECT 110.200 146.800 110.600 147.200 ;
        RECT 121.400 147.100 121.700 147.800 ;
        RECT 124.600 147.100 125.000 147.200 ;
        RECT 134.200 147.100 134.600 147.200 ;
        RECT 121.400 146.800 134.600 147.100 ;
        RECT 161.400 147.100 161.800 147.200 ;
        RECT 167.000 147.100 167.300 147.800 ;
        RECT 161.400 146.800 167.300 147.100 ;
        RECT 83.800 146.100 84.200 146.200 ;
        RECT 79.800 145.800 84.200 146.100 ;
        RECT 87.000 146.100 87.400 146.200 ;
        RECT 91.800 146.100 92.200 146.200 ;
        RECT 87.000 145.800 92.200 146.100 ;
        RECT 94.200 146.100 94.600 146.200 ;
        RECT 96.600 146.100 97.000 146.200 ;
        RECT 94.200 145.800 97.000 146.100 ;
        RECT 99.000 146.100 99.400 146.200 ;
        RECT 110.200 146.100 110.500 146.800 ;
        RECT 119.000 146.100 119.400 146.300 ;
        RECT 123.000 146.100 123.400 146.200 ;
        RECT 99.000 145.800 107.300 146.100 ;
        RECT 110.200 145.800 123.400 146.100 ;
        RECT 148.600 146.100 149.000 146.200 ;
        RECT 162.200 146.100 162.600 146.200 ;
        RECT 173.400 146.100 173.800 146.200 ;
        RECT 148.600 145.800 173.800 146.100 ;
        RECT 107.000 145.200 107.300 145.800 ;
        RECT 37.400 145.100 37.800 145.200 ;
        RECT 55.800 145.100 56.200 145.200 ;
        RECT 71.800 145.100 72.200 145.200 ;
        RECT 88.600 145.100 89.000 145.200 ;
        RECT 37.400 144.800 89.000 145.100 ;
        RECT 94.200 145.100 94.600 145.200 ;
        RECT 95.800 145.100 96.200 145.200 ;
        RECT 94.200 144.800 96.200 145.100 ;
        RECT 107.000 145.100 107.400 145.200 ;
        RECT 124.600 145.100 125.000 145.200 ;
        RECT 135.800 145.100 136.200 145.200 ;
        RECT 151.800 145.100 152.200 145.200 ;
        RECT 107.000 144.800 152.200 145.100 ;
        RECT 162.200 145.100 162.600 145.200 ;
        RECT 163.000 145.100 163.400 145.200 ;
        RECT 166.200 145.100 166.600 145.200 ;
        RECT 170.200 145.100 170.600 145.200 ;
        RECT 175.000 145.100 175.400 145.200 ;
        RECT 184.600 145.100 185.000 145.200 ;
        RECT 162.200 144.800 163.400 145.100 ;
        RECT 165.400 144.800 170.600 145.100 ;
        RECT 171.000 144.800 185.000 145.100 ;
        RECT 171.000 144.200 171.300 144.800 ;
        RECT 1.400 144.100 1.800 144.200 ;
        RECT 12.600 144.100 13.000 144.200 ;
        RECT 13.400 144.100 13.800 144.200 ;
        RECT 1.400 143.800 13.800 144.100 ;
        RECT 39.000 144.100 39.400 144.200 ;
        RECT 42.200 144.100 42.600 144.200 ;
        RECT 51.800 144.100 52.200 144.200 ;
        RECT 39.000 143.800 52.200 144.100 ;
        RECT 63.000 144.100 63.400 144.200 ;
        RECT 80.600 144.100 81.000 144.200 ;
        RECT 63.000 143.800 81.000 144.100 ;
        RECT 83.000 144.100 83.400 144.200 ;
        RECT 85.400 144.100 85.800 144.200 ;
        RECT 83.000 143.800 85.800 144.100 ;
        RECT 171.000 143.800 171.400 144.200 ;
        RECT 38.200 143.100 38.600 143.200 ;
        RECT 63.800 143.100 64.200 143.200 ;
        RECT 38.200 142.800 64.200 143.100 ;
        RECT 73.400 143.100 73.800 143.200 ;
        RECT 86.200 143.100 86.600 143.200 ;
        RECT 73.400 142.800 86.600 143.100 ;
        RECT 90.200 143.100 90.600 143.200 ;
        RECT 93.400 143.100 93.800 143.200 ;
        RECT 90.200 142.800 93.800 143.100 ;
        RECT 119.800 143.100 120.200 143.200 ;
        RECT 127.800 143.100 128.200 143.200 ;
        RECT 119.800 142.800 128.200 143.100 ;
        RECT 138.200 143.100 138.600 143.200 ;
        RECT 163.800 143.100 164.200 143.200 ;
        RECT 180.600 143.100 181.000 143.200 ;
        RECT 190.200 143.100 190.600 143.200 ;
        RECT 138.200 142.800 190.600 143.100 ;
        RECT 18.200 142.100 18.600 142.200 ;
        RECT 27.000 142.100 27.400 142.200 ;
        RECT 18.200 141.800 27.400 142.100 ;
        RECT 75.000 142.100 75.400 142.200 ;
        RECT 81.400 142.100 81.800 142.200 ;
        RECT 75.000 141.800 81.800 142.100 ;
        RECT 127.800 142.100 128.200 142.200 ;
        RECT 131.800 142.100 132.200 142.200 ;
        RECT 127.800 141.800 132.200 142.100 ;
        RECT 66.200 141.100 66.600 141.200 ;
        RECT 90.200 141.100 90.600 141.200 ;
        RECT 66.200 140.800 90.600 141.100 ;
        RECT 7.000 140.100 7.400 140.200 ;
        RECT 25.400 140.100 25.800 140.200 ;
        RECT 28.600 140.100 29.000 140.200 ;
        RECT 7.000 139.800 29.000 140.100 ;
        RECT 51.800 140.100 52.200 140.200 ;
        RECT 54.200 140.100 54.600 140.200 ;
        RECT 57.400 140.100 57.800 140.200 ;
        RECT 51.800 139.800 57.800 140.100 ;
        RECT 35.800 139.100 36.200 139.200 ;
        RECT 44.600 139.100 45.000 139.200 ;
        RECT 63.000 139.100 63.400 139.200 ;
        RECT 35.800 138.800 63.400 139.100 ;
        RECT 159.000 139.100 159.400 139.200 ;
        RECT 161.400 139.100 161.800 139.200 ;
        RECT 159.000 138.800 161.800 139.100 ;
        RECT 70.200 138.100 70.600 138.200 ;
        RECT 79.000 138.100 79.400 138.200 ;
        RECT 100.600 138.100 101.000 138.200 ;
        RECT 70.200 137.800 101.000 138.100 ;
        RECT 111.800 138.100 112.200 138.200 ;
        RECT 131.000 138.100 131.400 138.200 ;
        RECT 161.400 138.100 161.800 138.200 ;
        RECT 173.400 138.100 173.800 138.200 ;
        RECT 111.800 137.800 173.800 138.100 ;
        RECT 15.800 137.100 16.200 137.200 ;
        RECT 38.200 137.100 38.600 137.200 ;
        RECT 15.800 136.800 38.600 137.100 ;
        RECT 66.200 137.100 66.600 137.200 ;
        RECT 71.000 137.100 71.400 137.200 ;
        RECT 66.200 136.800 71.400 137.100 ;
        RECT 71.800 136.800 72.200 137.200 ;
        RECT 73.400 137.100 73.800 137.200 ;
        RECT 74.200 137.100 74.600 137.200 ;
        RECT 137.400 137.100 137.800 137.200 ;
        RECT 73.400 136.800 74.600 137.100 ;
        RECT 131.800 136.800 137.800 137.100 ;
        RECT 145.400 137.100 145.800 137.200 ;
        RECT 149.400 137.100 149.800 137.200 ;
        RECT 145.400 136.800 149.800 137.100 ;
        RECT 0.600 136.100 1.000 136.200 ;
        RECT 19.000 136.100 19.400 136.200 ;
        RECT 23.000 136.100 23.400 136.200 ;
        RECT 0.600 135.800 23.400 136.100 ;
        RECT 27.000 136.100 27.400 136.200 ;
        RECT 27.800 136.100 28.200 136.200 ;
        RECT 27.000 135.800 28.200 136.100 ;
        RECT 37.400 136.100 37.800 136.200 ;
        RECT 43.800 136.100 44.200 136.200 ;
        RECT 37.400 135.800 44.200 136.100 ;
        RECT 56.600 136.100 57.000 136.200 ;
        RECT 61.400 136.100 61.800 136.200 ;
        RECT 63.800 136.100 64.200 136.200 ;
        RECT 71.800 136.100 72.100 136.800 ;
        RECT 131.800 136.200 132.100 136.800 ;
        RECT 56.600 135.800 72.100 136.100 ;
        RECT 101.400 135.800 101.800 136.200 ;
        RECT 113.400 136.100 113.800 136.200 ;
        RECT 125.400 136.100 125.800 136.200 ;
        RECT 113.400 135.800 125.800 136.100 ;
        RECT 131.800 135.800 132.200 136.200 ;
        RECT 134.200 136.100 134.600 136.200 ;
        RECT 154.200 136.100 154.600 136.200 ;
        RECT 157.400 136.100 157.800 136.200 ;
        RECT 160.600 136.100 161.000 136.200 ;
        RECT 134.200 135.800 161.000 136.100 ;
        RECT 11.800 135.100 12.200 135.200 ;
        RECT 12.600 135.100 13.000 135.200 ;
        RECT 30.200 135.100 30.600 135.200 ;
        RECT 31.800 135.100 32.200 135.200 ;
        RECT 11.800 134.800 22.500 135.100 ;
        RECT 30.200 134.800 32.200 135.100 ;
        RECT 63.000 135.100 63.400 135.200 ;
        RECT 67.800 135.100 68.200 135.200 ;
        RECT 69.400 135.100 69.800 135.200 ;
        RECT 63.000 134.800 69.800 135.100 ;
        RECT 71.000 135.100 71.400 135.200 ;
        RECT 75.800 135.100 76.200 135.200 ;
        RECT 71.000 134.800 76.200 135.100 ;
        RECT 84.600 134.800 85.000 135.200 ;
        RECT 92.600 135.100 93.000 135.200 ;
        RECT 93.400 135.100 93.800 135.200 ;
        RECT 92.600 134.800 93.800 135.100 ;
        RECT 96.600 135.100 97.000 135.200 ;
        RECT 101.400 135.100 101.700 135.800 ;
        RECT 96.600 134.800 101.700 135.100 ;
        RECT 105.400 135.100 105.800 135.200 ;
        RECT 123.000 135.100 123.400 135.200 ;
        RECT 123.800 135.100 124.200 135.200 ;
        RECT 130.200 135.100 130.600 135.200 ;
        RECT 105.400 134.800 124.200 135.100 ;
        RECT 127.000 134.800 130.600 135.100 ;
        RECT 133.400 135.100 133.800 135.200 ;
        RECT 136.600 135.100 137.000 135.200 ;
        RECT 138.200 135.100 138.600 135.200 ;
        RECT 141.400 135.100 141.800 135.200 ;
        RECT 133.400 134.800 141.800 135.100 ;
        RECT 143.000 134.800 143.400 135.200 ;
        RECT 164.600 135.100 165.000 135.200 ;
        RECT 165.400 135.100 165.800 135.200 ;
        RECT 164.600 134.800 165.800 135.100 ;
        RECT 166.200 135.100 166.600 135.200 ;
        RECT 168.600 135.100 169.000 135.200 ;
        RECT 166.200 134.800 169.000 135.100 ;
        RECT 172.600 135.100 173.000 135.200 ;
        RECT 184.600 135.100 185.000 135.200 ;
        RECT 172.600 134.800 185.000 135.100 ;
        RECT 22.200 134.200 22.500 134.800 ;
        RECT 6.200 134.100 6.600 134.200 ;
        RECT 13.400 134.100 13.800 134.200 ;
        RECT 19.800 134.100 20.200 134.200 ;
        RECT 6.200 133.800 20.200 134.100 ;
        RECT 22.200 133.800 22.600 134.200 ;
        RECT 32.600 134.100 33.000 134.200 ;
        RECT 35.000 134.100 35.400 134.200 ;
        RECT 32.600 133.800 35.400 134.100 ;
        RECT 42.200 134.100 42.600 134.200 ;
        RECT 43.800 134.100 44.200 134.200 ;
        RECT 42.200 133.800 44.200 134.100 ;
        RECT 55.800 134.100 56.200 134.200 ;
        RECT 56.600 134.100 57.000 134.200 ;
        RECT 55.800 133.800 57.000 134.100 ;
        RECT 59.000 134.100 59.400 134.200 ;
        RECT 61.400 134.100 61.800 134.200 ;
        RECT 59.000 133.800 61.800 134.100 ;
        RECT 65.400 134.100 65.800 134.200 ;
        RECT 72.600 134.100 73.000 134.200 ;
        RECT 65.400 133.800 73.000 134.100 ;
        RECT 73.400 134.100 73.800 134.200 ;
        RECT 84.600 134.100 84.900 134.800 ;
        RECT 127.000 134.200 127.300 134.800 ;
        RECT 73.400 133.800 84.900 134.100 ;
        RECT 85.400 134.100 85.800 134.200 ;
        RECT 91.800 134.100 92.200 134.200 ;
        RECT 110.200 134.100 110.600 134.200 ;
        RECT 85.400 133.800 110.600 134.100 ;
        RECT 127.000 133.800 127.400 134.200 ;
        RECT 141.400 134.100 141.800 134.200 ;
        RECT 137.400 133.800 141.800 134.100 ;
        RECT 143.000 134.100 143.300 134.800 ;
        RECT 145.400 134.100 145.800 134.200 ;
        RECT 143.000 133.800 145.800 134.100 ;
        RECT 151.800 134.100 152.200 134.200 ;
        RECT 155.000 134.100 155.400 134.200 ;
        RECT 151.800 133.800 155.400 134.100 ;
        RECT 157.400 134.100 157.800 134.200 ;
        RECT 158.200 134.100 158.600 134.200 ;
        RECT 157.400 133.800 158.600 134.100 ;
        RECT 160.600 134.100 161.000 134.200 ;
        RECT 165.400 134.100 165.800 134.200 ;
        RECT 160.600 133.800 165.800 134.100 ;
        RECT 167.800 134.100 168.200 134.200 ;
        RECT 172.600 134.100 173.000 134.200 ;
        RECT 167.800 133.800 173.000 134.100 ;
        RECT 180.600 134.100 181.000 134.200 ;
        RECT 183.000 134.100 183.400 134.200 ;
        RECT 180.600 133.800 183.400 134.100 ;
        RECT 137.400 133.200 137.700 133.800 ;
        RECT 14.200 133.100 14.600 133.200 ;
        RECT 19.000 133.100 19.400 133.200 ;
        RECT 20.600 133.100 21.000 133.200 ;
        RECT 14.200 132.800 21.000 133.100 ;
        RECT 21.400 133.100 21.800 133.200 ;
        RECT 24.600 133.100 25.000 133.200 ;
        RECT 21.400 132.800 25.000 133.100 ;
        RECT 30.200 132.800 30.600 133.200 ;
        RECT 37.400 133.100 37.800 133.200 ;
        RECT 39.000 133.100 39.400 133.200 ;
        RECT 37.400 132.800 39.400 133.100 ;
        RECT 71.000 133.100 71.400 133.200 ;
        RECT 75.000 133.100 75.400 133.200 ;
        RECT 71.000 132.800 75.400 133.100 ;
        RECT 75.800 133.100 76.200 133.200 ;
        RECT 131.800 133.100 132.200 133.200 ;
        RECT 75.800 132.800 132.200 133.100 ;
        RECT 137.400 132.800 137.800 133.200 ;
        RECT 143.800 133.100 144.200 133.200 ;
        RECT 151.800 133.100 152.200 133.200 ;
        RECT 143.800 132.800 152.200 133.100 ;
        RECT 160.600 133.100 161.000 133.200 ;
        RECT 162.200 133.100 162.600 133.200 ;
        RECT 160.600 132.800 162.600 133.100 ;
        RECT 164.600 133.100 165.000 133.200 ;
        RECT 164.600 132.800 167.300 133.100 ;
        RECT 23.800 132.100 24.200 132.200 ;
        RECT 30.200 132.100 30.500 132.800 ;
        RECT 167.000 132.200 167.300 132.800 ;
        RECT 23.800 131.800 30.500 132.100 ;
        RECT 52.600 132.100 53.000 132.200 ;
        RECT 54.200 132.100 54.600 132.200 ;
        RECT 65.400 132.100 65.800 132.200 ;
        RECT 52.600 131.800 65.800 132.100 ;
        RECT 68.600 132.100 69.000 132.200 ;
        RECT 71.800 132.100 72.200 132.200 ;
        RECT 68.600 131.800 72.200 132.100 ;
        RECT 83.800 132.100 84.200 132.200 ;
        RECT 120.600 132.100 121.000 132.200 ;
        RECT 83.800 131.800 121.000 132.100 ;
        RECT 140.600 132.100 141.000 132.200 ;
        RECT 145.400 132.100 145.800 132.200 ;
        RECT 140.600 131.800 145.800 132.100 ;
        RECT 147.800 132.100 148.200 132.200 ;
        RECT 153.400 132.100 153.800 132.200 ;
        RECT 156.600 132.100 157.000 132.200 ;
        RECT 147.800 131.800 157.000 132.100 ;
        RECT 167.000 131.800 167.400 132.200 ;
        RECT 28.600 131.100 29.000 131.200 ;
        RECT 34.200 131.100 34.600 131.200 ;
        RECT 28.600 130.800 34.600 131.100 ;
        RECT 37.400 131.100 37.800 131.200 ;
        RECT 43.000 131.100 43.400 131.200 ;
        RECT 37.400 130.800 43.400 131.100 ;
        RECT 56.600 131.100 57.000 131.200 ;
        RECT 63.800 131.100 64.200 131.200 ;
        RECT 87.800 131.100 88.200 131.200 ;
        RECT 56.600 130.800 88.200 131.100 ;
        RECT 88.600 131.100 89.000 131.200 ;
        RECT 89.400 131.100 89.800 131.200 ;
        RECT 88.600 130.800 89.800 131.100 ;
        RECT 110.200 131.100 110.600 131.200 ;
        RECT 137.400 131.100 137.800 131.200 ;
        RECT 110.200 130.800 137.800 131.100 ;
        RECT 139.800 131.100 140.200 131.200 ;
        RECT 146.200 131.100 146.600 131.200 ;
        RECT 139.800 130.800 146.600 131.100 ;
        RECT 6.200 130.100 6.600 130.200 ;
        RECT 40.600 130.100 41.000 130.200 ;
        RECT 6.200 129.800 41.000 130.100 ;
        RECT 51.000 130.100 51.400 130.200 ;
        RECT 57.400 130.100 57.800 130.200 ;
        RECT 51.000 129.800 57.800 130.100 ;
        RECT 83.800 130.100 84.200 130.200 ;
        RECT 84.600 130.100 85.000 130.200 ;
        RECT 83.800 129.800 85.000 130.100 ;
        RECT 131.800 130.100 132.200 130.200 ;
        RECT 147.000 130.100 147.400 130.200 ;
        RECT 131.800 129.800 147.400 130.100 ;
        RECT 43.000 129.100 43.400 129.200 ;
        RECT 47.800 129.100 48.200 129.200 ;
        RECT 48.600 129.100 49.000 129.200 ;
        RECT 30.200 128.800 49.000 129.100 ;
        RECT 51.800 128.800 52.200 129.200 ;
        RECT 72.600 129.100 73.000 129.200 ;
        RECT 83.000 129.100 83.400 129.200 ;
        RECT 72.600 128.800 83.400 129.100 ;
        RECT 111.000 129.100 111.400 129.200 ;
        RECT 117.400 129.100 117.800 129.200 ;
        RECT 111.000 128.800 117.800 129.100 ;
        RECT 119.800 128.800 120.200 129.200 ;
        RECT 188.600 128.800 189.000 129.200 ;
        RECT 30.200 128.200 30.500 128.800 ;
        RECT 8.600 127.800 9.000 128.200 ;
        RECT 30.200 127.800 30.600 128.200 ;
        RECT 34.200 128.100 34.600 128.200 ;
        RECT 42.200 128.100 42.600 128.200 ;
        RECT 51.800 128.100 52.100 128.800 ;
        RECT 59.800 128.100 60.200 128.200 ;
        RECT 34.200 127.800 44.100 128.100 ;
        RECT 51.800 127.800 60.200 128.100 ;
        RECT 71.800 127.800 72.200 128.200 ;
        RECT 80.600 128.100 81.000 128.200 ;
        RECT 83.800 128.100 84.200 128.200 ;
        RECT 80.600 127.800 84.200 128.100 ;
        RECT 117.400 128.100 117.700 128.800 ;
        RECT 119.800 128.100 120.100 128.800 ;
        RECT 117.400 127.800 120.100 128.100 ;
        RECT 150.200 128.100 150.600 128.200 ;
        RECT 159.000 128.100 159.400 128.200 ;
        RECT 150.200 127.800 159.400 128.100 ;
        RECT 167.000 127.800 167.400 128.200 ;
        RECT 183.800 128.100 184.200 128.200 ;
        RECT 188.600 128.100 188.900 128.800 ;
        RECT 183.800 127.800 188.900 128.100 ;
        RECT 8.600 127.100 8.900 127.800 ;
        RECT 43.800 127.200 44.100 127.800 ;
        RECT 14.200 127.100 14.600 127.200 ;
        RECT 8.600 126.800 14.600 127.100 ;
        RECT 16.600 126.800 17.000 127.200 ;
        RECT 27.000 127.100 27.400 127.200 ;
        RECT 29.400 127.100 29.800 127.200 ;
        RECT 30.200 127.100 30.600 127.200 ;
        RECT 27.000 126.800 30.600 127.100 ;
        RECT 33.400 127.100 33.800 127.200 ;
        RECT 38.200 127.100 38.600 127.200 ;
        RECT 33.400 126.800 38.600 127.100 ;
        RECT 43.800 126.800 44.200 127.200 ;
        RECT 52.600 127.100 53.000 127.200 ;
        RECT 71.800 127.100 72.100 127.800 ;
        RECT 52.600 126.800 72.100 127.100 ;
        RECT 79.800 126.800 80.200 127.200 ;
        RECT 137.400 127.100 137.800 127.200 ;
        RECT 143.000 127.100 143.400 127.200 ;
        RECT 137.400 126.800 143.400 127.100 ;
        RECT 152.600 126.800 153.000 127.200 ;
        RECT 157.400 127.100 157.800 127.200 ;
        RECT 159.800 127.100 160.200 127.200 ;
        RECT 167.000 127.100 167.300 127.800 ;
        RECT 157.400 126.800 167.300 127.100 ;
        RECT 191.800 127.100 192.200 127.200 ;
        RECT 193.400 127.100 193.800 127.200 ;
        RECT 195.000 127.100 195.400 127.200 ;
        RECT 191.800 126.800 195.400 127.100 ;
        RECT 15.000 126.100 15.400 126.200 ;
        RECT 15.800 126.100 16.200 126.200 ;
        RECT 15.000 125.800 16.200 126.100 ;
        RECT 16.600 126.100 16.900 126.800 ;
        RECT 23.800 126.100 24.200 126.200 ;
        RECT 16.600 125.800 24.200 126.100 ;
        RECT 33.400 126.100 33.800 126.200 ;
        RECT 52.600 126.100 53.000 126.200 ;
        RECT 33.400 125.800 53.000 126.100 ;
        RECT 55.800 126.100 56.200 126.200 ;
        RECT 59.800 126.100 60.200 126.200 ;
        RECT 55.800 125.800 60.200 126.100 ;
        RECT 63.000 125.800 63.400 126.200 ;
        RECT 67.000 126.100 67.400 126.200 ;
        RECT 69.400 126.100 69.800 126.200 ;
        RECT 67.000 125.800 69.800 126.100 ;
        RECT 79.800 126.100 80.100 126.800 ;
        RECT 85.400 126.100 85.800 126.200 ;
        RECT 79.800 125.800 85.800 126.100 ;
        RECT 87.000 126.100 87.400 126.200 ;
        RECT 95.800 126.100 96.200 126.200 ;
        RECT 87.000 125.800 96.200 126.100 ;
        RECT 112.600 126.100 113.000 126.200 ;
        RECT 126.200 126.100 126.600 126.200 ;
        RECT 112.600 125.800 126.600 126.100 ;
        RECT 136.600 126.100 137.000 126.200 ;
        RECT 143.800 126.100 144.200 126.200 ;
        RECT 136.600 125.800 144.200 126.100 ;
        RECT 146.200 126.100 146.600 126.200 ;
        RECT 152.600 126.100 152.900 126.800 ;
        RECT 146.200 125.800 152.900 126.100 ;
        RECT 155.000 126.100 155.400 126.200 ;
        RECT 162.200 126.100 162.600 126.200 ;
        RECT 155.000 125.800 162.600 126.100 ;
        RECT 163.000 126.100 163.400 126.200 ;
        RECT 177.400 126.100 177.800 126.200 ;
        RECT 163.000 125.800 177.800 126.100 ;
        RECT 188.600 126.100 189.000 126.200 ;
        RECT 191.800 126.100 192.200 126.200 ;
        RECT 188.600 125.800 192.200 126.100 ;
        RECT 37.400 125.100 37.800 125.200 ;
        RECT 38.200 125.100 38.600 125.200 ;
        RECT 37.400 124.800 38.600 125.100 ;
        RECT 39.800 125.100 40.200 125.200 ;
        RECT 40.600 125.100 41.000 125.200 ;
        RECT 39.800 124.800 41.000 125.100 ;
        RECT 42.200 125.100 42.600 125.200 ;
        RECT 50.200 125.100 50.600 125.200 ;
        RECT 42.200 124.800 50.600 125.100 ;
        RECT 55.800 124.800 56.200 125.200 ;
        RECT 63.000 125.100 63.300 125.800 ;
        RECT 67.800 125.100 68.200 125.200 ;
        RECT 72.600 125.100 73.000 125.200 ;
        RECT 63.000 124.800 73.000 125.100 ;
        RECT 73.400 125.100 73.800 125.200 ;
        RECT 83.000 125.100 83.400 125.200 ;
        RECT 88.600 125.100 89.000 125.200 ;
        RECT 73.400 124.800 80.100 125.100 ;
        RECT 83.000 124.800 89.000 125.100 ;
        RECT 100.600 125.100 101.000 125.200 ;
        RECT 122.200 125.100 122.600 125.200 ;
        RECT 129.400 125.100 129.800 125.200 ;
        RECT 100.600 124.800 129.800 125.100 ;
        RECT 138.200 124.800 138.600 125.200 ;
        RECT 139.000 125.100 139.400 125.200 ;
        RECT 139.800 125.100 140.200 125.200 ;
        RECT 139.000 124.800 140.200 125.100 ;
        RECT 147.800 125.100 148.200 125.200 ;
        RECT 159.000 125.100 159.400 125.200 ;
        RECT 160.600 125.100 161.000 125.200 ;
        RECT 171.800 125.100 172.200 125.200 ;
        RECT 179.000 125.100 179.400 125.200 ;
        RECT 147.800 124.800 156.100 125.100 ;
        RECT 159.000 124.800 179.400 125.100 ;
        RECT 1.400 124.100 1.800 124.200 ;
        RECT 8.600 124.100 9.000 124.200 ;
        RECT 33.400 124.100 33.800 124.200 ;
        RECT 1.400 123.800 33.800 124.100 ;
        RECT 39.000 124.100 39.400 124.200 ;
        RECT 40.600 124.100 41.000 124.200 ;
        RECT 39.000 123.800 41.000 124.100 ;
        RECT 55.800 124.100 56.100 124.800 ;
        RECT 79.800 124.200 80.100 124.800 ;
        RECT 138.200 124.200 138.500 124.800 ;
        RECT 155.800 124.200 156.100 124.800 ;
        RECT 59.000 124.100 59.400 124.200 ;
        RECT 55.800 123.800 59.400 124.100 ;
        RECT 59.800 124.100 60.200 124.200 ;
        RECT 78.200 124.100 78.600 124.200 ;
        RECT 59.800 123.800 78.600 124.100 ;
        RECT 79.800 123.800 80.200 124.200 ;
        RECT 91.000 123.800 91.400 124.200 ;
        RECT 111.800 124.100 112.200 124.200 ;
        RECT 132.600 124.100 133.000 124.200 ;
        RECT 111.800 123.800 133.000 124.100 ;
        RECT 138.200 123.800 138.600 124.200 ;
        RECT 155.800 123.800 156.200 124.200 ;
        RECT 165.400 124.100 165.800 124.200 ;
        RECT 171.800 124.100 172.200 124.200 ;
        RECT 183.000 124.100 183.400 124.200 ;
        RECT 165.400 123.800 183.400 124.100 ;
        RECT 189.400 124.100 189.800 124.200 ;
        RECT 193.400 124.100 193.800 124.200 ;
        RECT 189.400 123.800 193.800 124.100 ;
        RECT 57.400 123.100 57.800 123.200 ;
        RECT 67.000 123.100 67.400 123.200 ;
        RECT 57.400 122.800 67.400 123.100 ;
        RECT 69.400 123.100 69.800 123.200 ;
        RECT 76.600 123.100 77.000 123.200 ;
        RECT 91.000 123.100 91.300 123.800 ;
        RECT 69.400 122.800 91.300 123.100 ;
        RECT 127.800 123.100 128.200 123.200 ;
        RECT 128.600 123.100 129.000 123.200 ;
        RECT 127.800 122.800 129.000 123.100 ;
        RECT 115.800 122.100 116.200 122.200 ;
        RECT 126.200 122.100 126.600 122.200 ;
        RECT 165.400 122.100 165.800 122.200 ;
        RECT 174.200 122.100 174.600 122.200 ;
        RECT 179.000 122.100 179.400 122.200 ;
        RECT 115.800 121.800 179.400 122.100 ;
        RECT 47.800 121.100 48.200 121.200 ;
        RECT 55.000 121.100 55.400 121.200 ;
        RECT 47.800 120.800 55.400 121.100 ;
        RECT 140.600 121.100 141.000 121.200 ;
        RECT 143.000 121.100 143.400 121.200 ;
        RECT 145.400 121.100 145.800 121.200 ;
        RECT 140.600 120.800 145.800 121.100 ;
        RECT 47.800 120.100 48.200 120.200 ;
        RECT 56.600 120.100 57.000 120.200 ;
        RECT 47.800 119.800 57.000 120.100 ;
        RECT 81.400 120.100 81.800 120.200 ;
        RECT 82.200 120.100 82.600 120.200 ;
        RECT 81.400 119.800 82.600 120.100 ;
        RECT 51.800 118.800 52.200 119.200 ;
        RECT 139.800 119.100 140.200 119.200 ;
        RECT 163.800 119.100 164.200 119.200 ;
        RECT 139.800 118.800 164.200 119.100 ;
        RECT 39.800 118.100 40.200 118.200 ;
        RECT 51.800 118.100 52.100 118.800 ;
        RECT 39.800 117.800 52.100 118.100 ;
        RECT 75.800 118.100 76.200 118.200 ;
        RECT 87.000 118.100 87.400 118.200 ;
        RECT 75.800 117.800 87.400 118.100 ;
        RECT 110.200 118.100 110.600 118.200 ;
        RECT 123.800 118.100 124.200 118.200 ;
        RECT 127.800 118.100 128.200 118.200 ;
        RECT 110.200 117.800 128.200 118.100 ;
        RECT 131.000 118.100 131.400 118.200 ;
        RECT 182.200 118.100 182.600 118.200 ;
        RECT 186.200 118.100 186.600 118.200 ;
        RECT 131.000 117.800 186.600 118.100 ;
        RECT 9.400 117.100 9.800 117.200 ;
        RECT 10.200 117.100 10.600 117.200 ;
        RECT 28.600 117.100 29.000 117.200 ;
        RECT 9.400 116.800 29.000 117.100 ;
        RECT 42.200 117.100 42.600 117.200 ;
        RECT 43.800 117.100 44.200 117.200 ;
        RECT 48.600 117.100 49.000 117.200 ;
        RECT 51.800 117.100 52.200 117.200 ;
        RECT 42.200 116.800 49.000 117.100 ;
        RECT 51.000 116.800 52.200 117.100 ;
        RECT 65.400 117.100 65.800 117.200 ;
        RECT 68.600 117.100 69.000 117.200 ;
        RECT 79.800 117.100 80.200 117.200 ;
        RECT 83.800 117.100 84.200 117.200 ;
        RECT 65.400 116.800 84.200 117.100 ;
        RECT 103.000 117.100 103.400 117.200 ;
        RECT 113.400 117.100 113.800 117.200 ;
        RECT 103.000 116.800 113.800 117.100 ;
        RECT 127.800 116.800 128.200 117.200 ;
        RECT 131.000 117.100 131.400 117.200 ;
        RECT 150.200 117.100 150.600 117.200 ;
        RECT 131.000 116.800 150.600 117.100 ;
        RECT 175.000 117.100 175.400 117.200 ;
        RECT 177.400 117.100 177.800 117.200 ;
        RECT 175.000 116.800 177.800 117.100 ;
        RECT 28.600 115.800 29.000 116.200 ;
        RECT 45.400 116.100 45.800 116.200 ;
        RECT 50.200 116.100 50.600 116.200 ;
        RECT 55.000 116.100 55.400 116.200 ;
        RECT 45.400 115.800 50.600 116.100 ;
        RECT 51.000 115.800 55.400 116.100 ;
        RECT 59.800 116.100 60.200 116.200 ;
        RECT 62.200 116.100 62.600 116.200 ;
        RECT 59.800 115.800 62.600 116.100 ;
        RECT 80.600 116.100 81.000 116.200 ;
        RECT 86.200 116.100 86.600 116.200 ;
        RECT 112.600 116.100 113.000 116.200 ;
        RECT 80.600 115.800 113.000 116.100 ;
        RECT 125.400 116.100 125.800 116.200 ;
        RECT 127.800 116.100 128.100 116.800 ;
        RECT 125.400 115.800 128.100 116.100 ;
        RECT 135.800 116.100 136.200 116.200 ;
        RECT 155.800 116.100 156.200 116.200 ;
        RECT 135.800 115.800 156.200 116.100 ;
        RECT 156.600 116.100 157.000 116.200 ;
        RECT 168.600 116.100 169.000 116.200 ;
        RECT 172.600 116.100 173.000 116.200 ;
        RECT 183.800 116.100 184.200 116.200 ;
        RECT 186.200 116.100 186.600 116.200 ;
        RECT 156.600 115.800 173.000 116.100 ;
        RECT 179.800 115.800 183.300 116.100 ;
        RECT 183.800 115.800 186.600 116.100 ;
        RECT 12.600 115.100 13.000 115.200 ;
        RECT 13.400 115.100 13.800 115.200 ;
        RECT 12.600 114.800 13.800 115.100 ;
        RECT 25.400 115.100 25.800 115.200 ;
        RECT 28.600 115.100 28.900 115.800 ;
        RECT 25.400 114.800 28.900 115.100 ;
        RECT 35.000 115.100 35.400 115.200 ;
        RECT 35.800 115.100 36.200 115.200 ;
        RECT 35.000 114.800 36.200 115.100 ;
        RECT 49.400 115.100 49.800 115.200 ;
        RECT 51.000 115.100 51.300 115.800 ;
        RECT 49.400 114.800 51.300 115.100 ;
        RECT 54.200 115.100 54.600 115.200 ;
        RECT 58.200 115.100 58.600 115.200 ;
        RECT 54.200 114.800 58.600 115.100 ;
        RECT 59.800 115.100 60.200 115.200 ;
        RECT 61.400 115.100 61.800 115.200 ;
        RECT 71.000 115.100 71.400 115.200 ;
        RECT 83.800 115.100 84.200 115.200 ;
        RECT 59.800 114.800 71.400 115.100 ;
        RECT 81.400 114.800 84.200 115.100 ;
        RECT 107.000 115.100 107.400 115.200 ;
        RECT 109.400 115.100 109.800 115.200 ;
        RECT 107.000 114.800 109.800 115.100 ;
        RECT 114.200 115.100 114.600 115.200 ;
        RECT 129.400 115.100 129.800 115.200 ;
        RECT 114.200 114.800 129.800 115.100 ;
        RECT 130.200 115.100 130.600 115.200 ;
        RECT 131.000 115.100 131.400 115.200 ;
        RECT 130.200 114.800 131.400 115.100 ;
        RECT 137.400 115.100 137.800 115.200 ;
        RECT 142.200 115.100 142.600 115.200 ;
        RECT 151.800 115.100 152.200 115.200 ;
        RECT 156.600 115.100 156.900 115.800 ;
        RECT 179.800 115.200 180.100 115.800 ;
        RECT 183.000 115.200 183.300 115.800 ;
        RECT 173.400 115.100 173.800 115.200 ;
        RECT 137.400 114.800 140.100 115.100 ;
        RECT 142.200 114.800 156.900 115.100 ;
        RECT 164.600 114.800 173.800 115.100 ;
        RECT 179.800 114.800 180.200 115.200 ;
        RECT 183.000 114.800 183.400 115.200 ;
        RECT 185.400 115.100 185.800 115.200 ;
        RECT 189.400 115.100 189.800 115.200 ;
        RECT 185.400 114.800 189.800 115.100 ;
        RECT 10.200 114.100 10.600 114.200 ;
        RECT 11.800 114.100 12.200 114.200 ;
        RECT 12.600 114.100 13.000 114.200 ;
        RECT 10.200 113.800 13.000 114.100 ;
        RECT 14.200 114.100 14.600 114.400 ;
        RECT 81.400 114.200 81.700 114.800 ;
        RECT 139.800 114.200 140.100 114.800 ;
        RECT 164.600 114.700 165.000 114.800 ;
        RECT 27.000 114.100 27.400 114.200 ;
        RECT 14.200 113.800 27.400 114.100 ;
        RECT 35.800 114.100 36.200 114.200 ;
        RECT 40.600 114.100 41.000 114.200 ;
        RECT 35.800 113.800 41.000 114.100 ;
        RECT 51.000 114.100 51.400 114.200 ;
        RECT 63.000 114.100 63.400 114.200 ;
        RECT 51.000 113.800 63.400 114.100 ;
        RECT 81.400 113.800 81.800 114.200 ;
        RECT 86.200 114.100 86.600 114.200 ;
        RECT 87.000 114.100 87.400 114.200 ;
        RECT 86.200 113.800 87.400 114.100 ;
        RECT 107.800 114.100 108.200 114.200 ;
        RECT 120.600 114.100 121.000 114.200 ;
        RECT 124.600 114.100 125.000 114.200 ;
        RECT 107.800 113.800 125.000 114.100 ;
        RECT 129.400 114.100 129.800 114.200 ;
        RECT 135.000 114.100 135.400 114.200 ;
        RECT 129.400 113.800 135.400 114.100 ;
        RECT 139.800 114.100 140.200 114.200 ;
        RECT 149.400 114.100 149.800 114.200 ;
        RECT 174.200 114.100 174.600 114.200 ;
        RECT 139.800 113.800 149.800 114.100 ;
        RECT 154.200 113.800 174.600 114.100 ;
        RECT 183.000 114.100 183.300 114.800 ;
        RECT 188.600 114.100 189.000 114.200 ;
        RECT 183.000 113.800 189.000 114.100 ;
        RECT 154.200 113.200 154.500 113.800 ;
        RECT 19.000 113.100 19.400 113.200 ;
        RECT 31.800 113.100 32.200 113.200 ;
        RECT 56.600 113.100 57.000 113.200 ;
        RECT 60.600 113.100 61.000 113.200 ;
        RECT 19.000 112.800 39.300 113.100 ;
        RECT 56.600 112.800 61.000 113.100 ;
        RECT 77.400 113.100 77.800 113.200 ;
        RECT 91.000 113.100 91.400 113.200 ;
        RECT 93.400 113.100 93.800 113.200 ;
        RECT 98.200 113.100 98.600 113.200 ;
        RECT 77.400 112.800 98.600 113.100 ;
        RECT 110.200 113.100 110.600 113.200 ;
        RECT 113.400 113.100 113.800 113.200 ;
        RECT 110.200 112.800 113.800 113.100 ;
        RECT 154.200 112.800 154.600 113.200 ;
        RECT 167.000 113.100 167.400 113.200 ;
        RECT 169.400 113.100 169.800 113.200 ;
        RECT 176.600 113.100 177.000 113.200 ;
        RECT 180.600 113.100 181.000 113.200 ;
        RECT 167.000 112.800 181.000 113.100 ;
        RECT 185.400 113.100 185.800 113.200 ;
        RECT 190.200 113.100 190.600 113.200 ;
        RECT 194.200 113.100 194.600 113.200 ;
        RECT 185.400 112.800 194.600 113.100 ;
        RECT 39.000 112.200 39.300 112.800 ;
        RECT 39.000 111.800 39.400 112.200 ;
        RECT 57.400 112.100 57.800 112.200 ;
        RECT 66.200 112.100 66.600 112.200 ;
        RECT 57.400 111.800 66.600 112.100 ;
        RECT 67.000 112.100 67.400 112.200 ;
        RECT 85.400 112.100 85.800 112.200 ;
        RECT 67.000 111.800 85.800 112.100 ;
        RECT 101.400 112.100 101.800 112.200 ;
        RECT 110.200 112.100 110.600 112.200 ;
        RECT 101.400 111.800 110.600 112.100 ;
        RECT 123.000 112.100 123.400 112.200 ;
        RECT 123.800 112.100 124.200 112.200 ;
        RECT 123.000 111.800 124.200 112.100 ;
        RECT 152.600 112.100 153.000 112.200 ;
        RECT 164.600 112.100 165.000 112.200 ;
        RECT 152.600 111.800 165.000 112.100 ;
        RECT 25.400 111.100 25.800 111.200 ;
        RECT 51.000 111.100 51.400 111.200 ;
        RECT 25.400 110.800 51.400 111.100 ;
        RECT 62.200 111.100 62.600 111.200 ;
        RECT 67.800 111.100 68.200 111.200 ;
        RECT 62.200 110.800 68.200 111.100 ;
        RECT 79.800 111.100 80.200 111.200 ;
        RECT 89.400 111.100 89.800 111.200 ;
        RECT 95.000 111.100 95.400 111.200 ;
        RECT 79.800 110.800 95.400 111.100 ;
        RECT 112.600 111.100 113.000 111.200 ;
        RECT 123.000 111.100 123.400 111.200 ;
        RECT 112.600 110.800 123.400 111.100 ;
        RECT 126.200 111.100 126.600 111.200 ;
        RECT 171.800 111.100 172.200 111.200 ;
        RECT 126.200 110.800 172.200 111.100 ;
        RECT 38.200 110.100 38.600 110.200 ;
        RECT 39.800 110.100 40.200 110.200 ;
        RECT 38.200 109.800 40.200 110.100 ;
        RECT 60.600 110.100 61.000 110.200 ;
        RECT 76.600 110.100 77.000 110.200 ;
        RECT 60.600 109.800 77.000 110.100 ;
        RECT 87.000 110.100 87.400 110.200 ;
        RECT 90.200 110.100 90.600 110.200 ;
        RECT 94.200 110.100 94.600 110.200 ;
        RECT 87.000 109.800 94.600 110.100 ;
        RECT 121.400 110.100 121.800 110.200 ;
        RECT 137.400 110.100 137.800 110.200 ;
        RECT 121.400 109.800 137.800 110.100 ;
        RECT 146.200 110.100 146.600 110.200 ;
        RECT 147.000 110.100 147.400 110.200 ;
        RECT 159.000 110.100 159.400 110.200 ;
        RECT 162.200 110.100 162.600 110.200 ;
        RECT 146.200 109.800 162.600 110.100 ;
        RECT 11.000 109.100 11.400 109.200 ;
        RECT 15.800 109.100 16.200 109.200 ;
        RECT 11.000 108.800 16.200 109.100 ;
        RECT 23.800 109.100 24.200 109.200 ;
        RECT 27.000 109.100 27.400 109.200 ;
        RECT 23.800 108.800 27.400 109.100 ;
        RECT 36.600 109.100 37.000 109.200 ;
        RECT 37.400 109.100 37.800 109.200 ;
        RECT 36.600 108.800 37.800 109.100 ;
        RECT 66.200 109.100 66.600 109.200 ;
        RECT 82.200 109.100 82.600 109.200 ;
        RECT 87.000 109.100 87.400 109.200 ;
        RECT 66.200 108.800 87.400 109.100 ;
        RECT 89.400 109.100 89.800 109.200 ;
        RECT 91.800 109.100 92.200 109.200 ;
        RECT 89.400 108.800 92.200 109.100 ;
        RECT 95.000 109.100 95.400 109.200 ;
        RECT 103.000 109.100 103.400 109.200 ;
        RECT 95.000 108.800 103.400 109.100 ;
        RECT 124.600 109.100 125.000 109.200 ;
        RECT 133.400 109.100 133.800 109.200 ;
        RECT 135.800 109.100 136.200 109.200 ;
        RECT 142.200 109.100 142.600 109.200 ;
        RECT 145.400 109.100 145.800 109.200 ;
        RECT 124.600 108.800 145.800 109.100 ;
        RECT 155.000 108.800 155.400 109.200 ;
        RECT 191.800 109.100 192.200 109.200 ;
        RECT 194.200 109.100 194.600 109.200 ;
        RECT 191.800 108.800 194.600 109.100 ;
        RECT 7.800 108.100 8.200 108.200 ;
        RECT 8.600 108.100 9.000 108.200 ;
        RECT 12.600 108.100 13.000 108.200 ;
        RECT 7.800 107.800 13.000 108.100 ;
        RECT 15.000 108.100 15.400 108.200 ;
        RECT 16.600 108.100 17.000 108.200 ;
        RECT 15.000 107.800 17.000 108.100 ;
        RECT 17.400 107.800 17.800 108.200 ;
        RECT 29.400 108.100 29.800 108.200 ;
        RECT 37.400 108.100 37.800 108.200 ;
        RECT 39.800 108.100 40.200 108.200 ;
        RECT 40.600 108.100 41.000 108.200 ;
        RECT 29.400 107.800 41.000 108.100 ;
        RECT 61.400 108.100 61.800 108.200 ;
        RECT 63.800 108.100 64.200 108.200 ;
        RECT 61.400 107.800 64.200 108.100 ;
        RECT 64.600 108.100 65.000 108.200 ;
        RECT 70.200 108.100 70.600 108.200 ;
        RECT 64.600 107.800 70.600 108.100 ;
        RECT 77.400 108.100 77.800 108.200 ;
        RECT 92.600 108.100 93.000 108.200 ;
        RECT 77.400 107.800 93.000 108.100 ;
        RECT 102.200 107.800 102.600 108.200 ;
        RECT 138.200 107.800 138.600 108.200 ;
        RECT 155.000 108.100 155.300 108.800 ;
        RECT 160.600 108.100 161.000 108.200 ;
        RECT 155.000 107.800 161.000 108.100 ;
        RECT 163.000 108.100 163.400 108.200 ;
        RECT 167.000 108.100 167.400 108.200 ;
        RECT 163.000 107.800 167.400 108.100 ;
        RECT 1.400 107.100 1.800 107.200 ;
        RECT 7.800 107.100 8.200 107.200 ;
        RECT 11.000 107.100 11.400 107.200 ;
        RECT 1.400 106.800 11.400 107.100 ;
        RECT 12.600 107.100 13.000 107.200 ;
        RECT 17.400 107.100 17.700 107.800 ;
        RECT 12.600 106.800 17.700 107.100 ;
        RECT 23.800 107.100 24.200 107.200 ;
        RECT 36.600 107.100 37.000 107.200 ;
        RECT 37.400 107.100 37.800 107.200 ;
        RECT 23.800 106.800 30.500 107.100 ;
        RECT 36.600 106.800 37.800 107.100 ;
        RECT 41.400 107.100 41.800 107.200 ;
        RECT 43.000 107.100 43.400 107.200 ;
        RECT 41.400 106.800 43.400 107.100 ;
        RECT 50.200 107.100 50.600 107.200 ;
        RECT 55.000 107.100 55.400 107.200 ;
        RECT 65.400 107.100 65.800 107.200 ;
        RECT 67.000 107.100 67.400 107.200 ;
        RECT 50.200 106.800 67.400 107.100 ;
        RECT 102.200 107.100 102.500 107.800 ;
        RECT 116.600 107.100 117.000 107.200 ;
        RECT 102.200 106.800 117.000 107.100 ;
        RECT 135.000 107.100 135.400 107.200 ;
        RECT 138.200 107.100 138.500 107.800 ;
        RECT 135.000 106.800 138.500 107.100 ;
        RECT 152.600 106.800 153.000 107.200 ;
        RECT 162.200 107.100 162.600 107.200 ;
        RECT 164.600 107.100 165.000 107.200 ;
        RECT 162.200 106.800 165.000 107.100 ;
        RECT 167.800 107.100 168.200 107.200 ;
        RECT 168.600 107.100 169.000 107.200 ;
        RECT 167.800 106.800 169.000 107.100 ;
        RECT 190.200 106.800 190.600 107.200 ;
        RECT 30.200 106.200 30.500 106.800 ;
        RECT 59.000 106.200 59.300 106.800 ;
        RECT 10.200 106.100 10.600 106.200 ;
        RECT 13.400 106.100 13.800 106.200 ;
        RECT 10.200 105.800 13.800 106.100 ;
        RECT 30.200 105.800 30.600 106.200 ;
        RECT 31.800 106.100 32.200 106.200 ;
        RECT 35.000 106.100 35.400 106.200 ;
        RECT 31.800 105.800 35.400 106.100 ;
        RECT 47.800 106.100 48.200 106.200 ;
        RECT 48.600 106.100 49.000 106.200 ;
        RECT 47.800 105.800 49.000 106.100 ;
        RECT 59.000 105.800 59.400 106.200 ;
        RECT 64.600 106.100 65.000 106.200 ;
        RECT 66.200 106.100 66.600 106.200 ;
        RECT 64.600 105.800 66.600 106.100 ;
        RECT 67.800 106.100 68.200 106.200 ;
        RECT 68.600 106.100 69.000 106.200 ;
        RECT 75.000 106.100 75.400 106.200 ;
        RECT 67.800 105.800 75.400 106.100 ;
        RECT 81.400 106.100 81.800 106.200 ;
        RECT 83.800 106.100 84.200 106.200 ;
        RECT 81.400 105.800 84.200 106.100 ;
        RECT 89.400 106.100 89.800 106.200 ;
        RECT 99.000 106.100 99.400 106.200 ;
        RECT 113.400 106.100 113.800 106.200 ;
        RECT 89.400 105.800 99.400 106.100 ;
        RECT 110.200 105.800 113.800 106.100 ;
        RECT 130.200 106.100 130.600 106.200 ;
        RECT 141.400 106.100 141.800 106.200 ;
        RECT 130.200 105.800 141.800 106.100 ;
        RECT 149.400 106.100 149.800 106.200 ;
        RECT 152.600 106.100 152.900 106.800 ;
        RECT 190.200 106.200 190.500 106.800 ;
        RECT 149.400 105.800 152.900 106.100 ;
        RECT 156.600 106.100 157.000 106.200 ;
        RECT 158.200 106.100 158.600 106.200 ;
        RECT 156.600 105.800 158.600 106.100 ;
        RECT 160.600 106.100 161.000 106.200 ;
        RECT 163.000 106.100 163.400 106.200 ;
        RECT 165.400 106.100 165.800 106.200 ;
        RECT 160.600 105.800 165.800 106.100 ;
        RECT 173.400 106.100 173.800 106.200 ;
        RECT 182.200 106.100 182.600 106.200 ;
        RECT 173.400 105.800 182.600 106.100 ;
        RECT 190.200 105.800 190.600 106.200 ;
        RECT 110.200 105.200 110.500 105.800 ;
        RECT 12.600 105.100 13.000 105.200 ;
        RECT 14.200 105.100 14.600 105.200 ;
        RECT 12.600 104.800 14.600 105.100 ;
        RECT 19.800 105.100 20.200 105.200 ;
        RECT 22.200 105.100 22.600 105.200 ;
        RECT 40.600 105.100 41.000 105.200 ;
        RECT 19.800 104.800 22.600 105.100 ;
        RECT 39.000 104.800 41.000 105.100 ;
        RECT 59.800 105.100 60.200 105.200 ;
        RECT 70.200 105.100 70.600 105.200 ;
        RECT 59.800 104.800 70.600 105.100 ;
        RECT 110.200 104.800 110.600 105.200 ;
        RECT 39.000 104.200 39.300 104.800 ;
        RECT 2.200 104.100 2.600 104.200 ;
        RECT 5.400 104.100 5.800 104.200 ;
        RECT 19.000 104.100 19.400 104.200 ;
        RECT 2.200 103.800 19.400 104.100 ;
        RECT 39.000 103.800 39.400 104.200 ;
        RECT 42.200 104.100 42.600 104.200 ;
        RECT 46.200 104.100 46.600 104.200 ;
        RECT 42.200 103.800 46.600 104.100 ;
        RECT 60.600 104.100 61.000 104.200 ;
        RECT 73.400 104.100 73.800 104.200 ;
        RECT 60.600 103.800 73.800 104.100 ;
        RECT 104.600 104.100 105.000 104.200 ;
        RECT 107.000 104.100 107.400 104.200 ;
        RECT 104.600 103.800 107.400 104.100 ;
        RECT 35.800 103.100 36.200 103.200 ;
        RECT 77.400 103.100 77.800 103.200 ;
        RECT 35.800 102.800 77.800 103.100 ;
        RECT 15.000 102.100 15.400 102.200 ;
        RECT 26.200 102.100 26.600 102.200 ;
        RECT 15.000 101.800 26.600 102.100 ;
        RECT 53.400 102.100 53.800 102.200 ;
        RECT 55.800 102.100 56.200 102.200 ;
        RECT 103.000 102.100 103.400 102.200 ;
        RECT 53.400 101.800 103.400 102.100 ;
        RECT 151.000 102.100 151.400 102.200 ;
        RECT 154.200 102.100 154.600 102.200 ;
        RECT 151.000 101.800 154.600 102.100 ;
        RECT 54.200 101.100 54.600 101.200 ;
        RECT 73.400 101.100 73.800 101.200 ;
        RECT 54.200 100.800 73.800 101.100 ;
        RECT 14.200 99.100 14.600 99.200 ;
        RECT 39.800 99.100 40.200 99.200 ;
        RECT 14.200 98.800 40.200 99.100 ;
        RECT 103.000 99.100 103.400 99.200 ;
        RECT 111.800 99.100 112.200 99.200 ;
        RECT 103.000 98.800 112.200 99.100 ;
        RECT 118.200 99.100 118.600 99.200 ;
        RECT 128.600 99.100 129.000 99.200 ;
        RECT 118.200 98.800 129.000 99.100 ;
        RECT 143.000 99.100 143.400 99.200 ;
        RECT 153.400 99.100 153.800 99.200 ;
        RECT 143.000 98.800 153.800 99.100 ;
        RECT 180.600 99.100 181.000 99.200 ;
        RECT 183.800 99.100 184.200 99.200 ;
        RECT 180.600 98.800 184.200 99.100 ;
        RECT 31.800 98.100 32.200 98.200 ;
        RECT 54.200 98.100 54.600 98.200 ;
        RECT 56.600 98.100 57.000 98.200 ;
        RECT 60.600 98.100 61.000 98.200 ;
        RECT 31.800 97.800 61.000 98.100 ;
        RECT 81.400 98.100 81.800 98.200 ;
        RECT 87.000 98.100 87.400 98.200 ;
        RECT 81.400 97.800 87.400 98.100 ;
        RECT 111.800 98.100 112.200 98.200 ;
        RECT 112.600 98.100 113.000 98.200 ;
        RECT 111.800 97.800 113.000 98.100 ;
        RECT 115.800 98.100 116.200 98.200 ;
        RECT 119.800 98.100 120.200 98.200 ;
        RECT 115.800 97.800 120.200 98.100 ;
        RECT 35.000 96.800 35.400 97.200 ;
        RECT 35.800 97.100 36.200 97.200 ;
        RECT 42.200 97.100 42.600 97.200 ;
        RECT 35.800 96.800 42.600 97.100 ;
        RECT 43.800 97.100 44.200 97.200 ;
        RECT 44.600 97.100 45.000 97.200 ;
        RECT 53.400 97.100 53.800 97.200 ;
        RECT 131.800 97.100 132.200 97.200 ;
        RECT 43.800 96.800 132.200 97.100 ;
        RECT 133.400 97.100 133.800 97.200 ;
        RECT 159.000 97.100 159.400 97.200 ;
        RECT 133.400 96.800 159.400 97.100 ;
        RECT 1.400 96.100 1.800 96.200 ;
        RECT 2.200 96.100 2.600 96.200 ;
        RECT 1.400 95.800 2.600 96.100 ;
        RECT 10.200 96.100 10.600 96.200 ;
        RECT 33.400 96.100 33.800 96.200 ;
        RECT 10.200 95.800 33.800 96.100 ;
        RECT 35.000 96.100 35.300 96.800 ;
        RECT 38.200 96.100 38.600 96.200 ;
        RECT 35.000 95.800 38.600 96.100 ;
        RECT 40.600 96.100 41.000 96.200 ;
        RECT 55.800 96.100 56.200 96.200 ;
        RECT 40.600 95.800 56.200 96.100 ;
        RECT 73.400 96.100 73.800 96.200 ;
        RECT 80.600 96.100 81.000 96.200 ;
        RECT 130.200 96.100 130.600 96.200 ;
        RECT 73.400 95.800 130.600 96.100 ;
        RECT 149.400 95.800 149.800 96.200 ;
        RECT 176.600 95.800 177.000 96.200 ;
        RECT 2.200 95.100 2.600 95.200 ;
        RECT 17.400 95.100 17.800 95.200 ;
        RECT 27.800 95.100 28.200 95.200 ;
        RECT 2.200 94.800 17.800 95.100 ;
        RECT 19.000 94.800 28.200 95.100 ;
        RECT 31.000 95.100 31.400 95.200 ;
        RECT 37.400 95.100 37.800 95.200 ;
        RECT 31.000 94.800 37.800 95.100 ;
        RECT 39.000 95.100 39.400 95.200 ;
        RECT 39.800 95.100 40.200 95.200 ;
        RECT 39.000 94.800 40.200 95.100 ;
        RECT 41.400 94.800 41.800 95.200 ;
        RECT 42.200 95.100 42.600 95.200 ;
        RECT 47.000 95.100 47.400 95.200 ;
        RECT 51.800 95.100 52.200 95.200 ;
        RECT 42.200 94.800 52.200 95.100 ;
        RECT 58.200 94.800 58.600 95.200 ;
        RECT 59.800 95.100 60.200 95.200 ;
        RECT 62.200 95.100 62.600 95.200 ;
        RECT 59.800 94.800 62.600 95.100 ;
        RECT 67.800 95.100 68.200 95.200 ;
        RECT 74.200 95.100 74.600 95.200 ;
        RECT 67.800 94.800 74.600 95.100 ;
        RECT 84.600 95.100 85.000 95.200 ;
        RECT 121.400 95.100 121.800 95.200 ;
        RECT 84.600 94.800 121.800 95.100 ;
        RECT 125.400 95.100 125.800 95.200 ;
        RECT 126.200 95.100 126.600 95.200 ;
        RECT 125.400 94.800 126.600 95.100 ;
        RECT 149.400 95.100 149.700 95.800 ;
        RECT 159.800 95.100 160.200 95.200 ;
        RECT 149.400 94.800 160.200 95.100 ;
        RECT 166.200 94.800 166.600 95.200 ;
        RECT 174.200 95.100 174.600 95.200 ;
        RECT 176.600 95.100 176.900 95.800 ;
        RECT 174.200 94.800 176.900 95.100 ;
        RECT 179.000 95.100 179.400 95.200 ;
        RECT 179.000 94.800 186.600 95.100 ;
        RECT 19.000 94.700 19.400 94.800 ;
        RECT 41.400 94.200 41.700 94.800 ;
        RECT 58.200 94.200 58.500 94.800 ;
        RECT 166.200 94.200 166.500 94.800 ;
        RECT 186.200 94.700 186.600 94.800 ;
        RECT 7.800 94.100 8.200 94.200 ;
        RECT 8.600 94.100 9.000 94.200 ;
        RECT 7.800 93.800 9.000 94.100 ;
        RECT 25.400 94.100 25.800 94.200 ;
        RECT 26.200 94.100 26.600 94.200 ;
        RECT 25.400 93.800 26.600 94.100 ;
        RECT 33.400 94.100 33.800 94.200 ;
        RECT 35.800 94.100 36.200 94.200 ;
        RECT 33.400 93.800 36.200 94.100 ;
        RECT 38.200 94.100 38.600 94.200 ;
        RECT 39.800 94.100 40.200 94.200 ;
        RECT 38.200 93.800 40.200 94.100 ;
        RECT 41.400 93.800 41.800 94.200 ;
        RECT 43.000 94.100 43.400 94.200 ;
        RECT 45.400 94.100 45.800 94.200 ;
        RECT 47.800 94.100 48.200 94.200 ;
        RECT 43.000 93.800 45.800 94.100 ;
        RECT 46.200 93.800 48.200 94.100 ;
        RECT 58.200 93.800 58.600 94.200 ;
        RECT 68.600 93.800 69.000 94.200 ;
        RECT 87.000 94.100 87.400 94.200 ;
        RECT 93.400 94.100 93.800 94.200 ;
        RECT 87.000 93.800 93.800 94.100 ;
        RECT 107.800 94.100 108.200 94.200 ;
        RECT 110.200 94.100 110.600 94.200 ;
        RECT 107.800 93.800 110.600 94.100 ;
        RECT 113.400 94.100 113.800 94.200 ;
        RECT 117.400 94.100 117.800 94.200 ;
        RECT 113.400 93.800 117.800 94.100 ;
        RECT 119.800 93.800 120.200 94.200 ;
        RECT 128.600 94.100 129.000 94.200 ;
        RECT 131.000 94.100 131.400 94.200 ;
        RECT 128.600 93.800 131.400 94.100 ;
        RECT 143.000 93.800 143.400 94.200 ;
        RECT 166.200 93.800 166.600 94.200 ;
        RECT 169.400 94.100 169.800 94.200 ;
        RECT 172.600 94.100 173.000 94.200 ;
        RECT 169.400 93.800 173.000 94.100 ;
        RECT 46.200 93.200 46.500 93.800 ;
        RECT 7.800 93.100 8.200 93.200 ;
        RECT 12.600 93.100 13.000 93.200 ;
        RECT 7.800 92.800 13.000 93.100 ;
        RECT 30.200 93.100 30.600 93.200 ;
        RECT 34.200 93.100 34.600 93.200 ;
        RECT 30.200 92.800 34.600 93.100 ;
        RECT 39.000 93.100 39.400 93.200 ;
        RECT 43.000 93.100 43.400 93.200 ;
        RECT 39.000 92.800 43.400 93.100 ;
        RECT 46.200 92.800 46.600 93.200 ;
        RECT 59.000 93.100 59.400 93.200 ;
        RECT 61.400 93.100 61.800 93.200 ;
        RECT 59.000 92.800 61.800 93.100 ;
        RECT 63.000 93.100 63.400 93.200 ;
        RECT 68.600 93.100 68.900 93.800 ;
        RECT 63.000 92.800 68.900 93.100 ;
        RECT 80.600 93.100 81.000 93.200 ;
        RECT 87.800 93.100 88.200 93.200 ;
        RECT 91.000 93.100 91.400 93.200 ;
        RECT 105.400 93.100 105.800 93.200 ;
        RECT 80.600 92.800 105.800 93.100 ;
        RECT 119.800 93.100 120.100 93.800 ;
        RECT 125.400 93.100 125.800 93.200 ;
        RECT 143.000 93.100 143.300 93.800 ;
        RECT 119.800 92.800 143.300 93.100 ;
        RECT 7.800 92.100 8.200 92.200 ;
        RECT 8.600 92.100 9.000 92.200 ;
        RECT 7.800 91.800 9.000 92.100 ;
        RECT 10.200 92.100 10.600 92.200 ;
        RECT 27.000 92.100 27.400 92.200 ;
        RECT 10.200 91.800 27.400 92.100 ;
        RECT 34.200 92.100 34.600 92.200 ;
        RECT 42.200 92.100 42.600 92.200 ;
        RECT 34.200 91.800 42.600 92.100 ;
        RECT 48.600 92.100 49.000 92.200 ;
        RECT 55.800 92.100 56.200 92.200 ;
        RECT 81.400 92.100 81.800 92.200 ;
        RECT 48.600 91.800 81.800 92.100 ;
        RECT 115.000 92.100 115.400 92.200 ;
        RECT 119.800 92.100 120.200 92.200 ;
        RECT 115.000 91.800 120.200 92.100 ;
        RECT 127.800 92.100 128.200 92.200 ;
        RECT 131.000 92.100 131.400 92.200 ;
        RECT 127.800 91.800 131.400 92.100 ;
        RECT 131.800 92.100 132.200 92.200 ;
        RECT 132.600 92.100 133.000 92.200 ;
        RECT 131.800 91.800 133.000 92.100 ;
        RECT 133.400 92.100 133.800 92.200 ;
        RECT 139.800 92.100 140.200 92.200 ;
        RECT 133.400 91.800 140.200 92.100 ;
        RECT 171.800 92.100 172.200 92.200 ;
        RECT 172.600 92.100 173.000 92.200 ;
        RECT 191.000 92.100 191.400 92.200 ;
        RECT 171.800 91.800 191.400 92.100 ;
        RECT 3.800 91.100 4.200 91.200 ;
        RECT 10.200 91.100 10.600 91.200 ;
        RECT 3.800 90.800 10.600 91.100 ;
        RECT 11.800 91.100 12.200 91.200 ;
        RECT 15.800 91.100 16.200 91.200 ;
        RECT 11.800 90.800 16.200 91.100 ;
        RECT 27.000 91.100 27.400 91.200 ;
        RECT 31.800 91.100 32.200 91.200 ;
        RECT 27.000 90.800 32.200 91.100 ;
        RECT 45.400 91.100 45.800 91.200 ;
        RECT 58.200 91.100 58.600 91.200 ;
        RECT 45.400 90.800 58.600 91.100 ;
        RECT 130.200 91.100 130.600 91.200 ;
        RECT 143.000 91.100 143.400 91.200 ;
        RECT 167.800 91.100 168.200 91.200 ;
        RECT 130.200 90.800 168.200 91.100 ;
        RECT 191.800 91.100 192.200 91.200 ;
        RECT 195.000 91.100 195.400 91.200 ;
        RECT 191.800 90.800 195.400 91.100 ;
        RECT 2.200 90.100 2.600 90.200 ;
        RECT 5.400 90.100 5.800 90.200 ;
        RECT 2.200 89.800 5.800 90.100 ;
        RECT 13.400 90.100 13.800 90.200 ;
        RECT 36.600 90.100 37.000 90.200 ;
        RECT 39.800 90.100 40.200 90.200 ;
        RECT 13.400 89.800 40.200 90.100 ;
        RECT 40.600 90.100 41.000 90.200 ;
        RECT 51.000 90.100 51.400 90.200 ;
        RECT 40.600 89.800 51.400 90.100 ;
        RECT 51.800 90.100 52.200 90.200 ;
        RECT 57.400 90.100 57.800 90.200 ;
        RECT 51.800 89.800 57.800 90.100 ;
        RECT 159.800 89.800 160.200 90.200 ;
        RECT 159.800 89.200 160.100 89.800 ;
        RECT 37.400 89.100 37.800 89.200 ;
        RECT 44.600 89.100 45.000 89.200 ;
        RECT 57.400 89.100 57.800 89.200 ;
        RECT 37.400 88.800 45.000 89.100 ;
        RECT 45.400 88.800 57.800 89.100 ;
        RECT 58.200 88.800 58.600 89.200 ;
        RECT 63.000 89.100 63.400 89.200 ;
        RECT 67.800 89.100 68.200 89.200 ;
        RECT 63.000 88.800 68.200 89.100 ;
        RECT 104.600 89.100 105.000 89.200 ;
        RECT 107.000 89.100 107.400 89.200 ;
        RECT 113.400 89.100 113.800 89.200 ;
        RECT 104.600 88.800 113.800 89.100 ;
        RECT 114.200 89.100 114.600 89.200 ;
        RECT 123.800 89.100 124.200 89.200 ;
        RECT 114.200 88.800 124.200 89.100 ;
        RECT 159.800 88.800 160.200 89.200 ;
        RECT 183.800 89.100 184.200 89.200 ;
        RECT 184.600 89.100 185.000 89.200 ;
        RECT 183.800 88.800 185.000 89.100 ;
        RECT 45.400 88.200 45.700 88.800 ;
        RECT 58.200 88.200 58.500 88.800 ;
        RECT 32.600 88.100 33.000 88.200 ;
        RECT 35.000 88.100 35.400 88.200 ;
        RECT 32.600 87.800 35.400 88.100 ;
        RECT 38.200 88.100 38.600 88.200 ;
        RECT 43.800 88.100 44.200 88.200 ;
        RECT 38.200 87.800 44.200 88.100 ;
        RECT 45.400 87.800 45.800 88.200 ;
        RECT 53.400 88.100 53.800 88.200 ;
        RECT 58.200 88.100 58.600 88.200 ;
        RECT 53.400 87.800 58.600 88.100 ;
        RECT 95.000 87.800 95.400 88.200 ;
        RECT 106.200 88.100 106.600 88.200 ;
        RECT 117.400 88.100 117.800 88.200 ;
        RECT 106.200 87.800 117.800 88.100 ;
        RECT 121.400 88.100 121.800 88.200 ;
        RECT 127.000 88.100 127.400 88.200 ;
        RECT 137.400 88.100 137.800 88.200 ;
        RECT 142.200 88.100 142.600 88.200 ;
        RECT 145.400 88.100 145.800 88.200 ;
        RECT 121.400 87.800 145.800 88.100 ;
        RECT 174.200 88.100 174.600 88.200 ;
        RECT 175.800 88.100 176.200 88.200 ;
        RECT 181.400 88.100 181.800 88.200 ;
        RECT 174.200 87.800 181.800 88.100 ;
        RECT 1.400 87.100 1.800 87.200 ;
        RECT 6.200 87.100 6.600 87.200 ;
        RECT 1.400 86.800 6.600 87.100 ;
        RECT 23.800 87.100 24.200 87.200 ;
        RECT 28.600 87.100 29.000 87.200 ;
        RECT 35.800 87.100 36.200 87.200 ;
        RECT 23.800 86.800 36.200 87.100 ;
        RECT 43.800 87.100 44.200 87.200 ;
        RECT 44.600 87.100 45.000 87.200 ;
        RECT 47.800 87.100 48.200 87.200 ;
        RECT 43.800 86.800 48.200 87.100 ;
        RECT 68.600 86.800 69.000 87.200 ;
        RECT 95.000 87.100 95.300 87.800 ;
        RECT 104.600 87.100 105.000 87.200 ;
        RECT 111.000 87.100 111.400 87.200 ;
        RECT 95.000 86.800 111.400 87.100 ;
        RECT 119.000 87.100 119.400 87.200 ;
        RECT 123.800 87.100 124.200 87.200 ;
        RECT 119.000 86.800 124.200 87.100 ;
        RECT 132.600 87.100 133.000 87.200 ;
        RECT 137.400 87.100 137.800 87.200 ;
        RECT 150.200 87.100 150.600 87.200 ;
        RECT 132.600 86.800 150.600 87.100 ;
        RECT 153.400 87.100 153.800 87.200 ;
        RECT 163.800 87.100 164.200 87.200 ;
        RECT 169.400 87.100 169.800 87.200 ;
        RECT 153.400 86.800 157.700 87.100 ;
        RECT 163.800 86.800 169.800 87.100 ;
        RECT 8.600 86.100 9.000 86.200 ;
        RECT 11.800 86.100 12.200 86.200 ;
        RECT 7.800 85.800 12.200 86.100 ;
        RECT 30.200 86.100 30.600 86.200 ;
        RECT 42.200 86.100 42.600 86.200 ;
        RECT 47.000 86.100 47.400 86.200 ;
        RECT 30.200 85.800 47.400 86.100 ;
        RECT 59.800 86.100 60.200 86.200 ;
        RECT 60.600 86.100 61.000 86.200 ;
        RECT 66.200 86.100 66.600 86.200 ;
        RECT 59.800 85.800 66.600 86.100 ;
        RECT 68.600 86.100 68.900 86.800 ;
        RECT 157.400 86.200 157.700 86.800 ;
        RECT 79.000 86.100 79.400 86.200 ;
        RECT 68.600 85.800 79.400 86.100 ;
        RECT 104.600 85.800 105.000 86.200 ;
        RECT 108.600 86.100 109.000 86.200 ;
        RECT 121.400 86.100 121.800 86.200 ;
        RECT 108.600 85.800 121.800 86.100 ;
        RECT 126.200 86.100 126.600 86.200 ;
        RECT 138.200 86.100 138.600 86.200 ;
        RECT 139.000 86.100 139.400 86.200 ;
        RECT 126.200 85.800 139.400 86.100 ;
        RECT 140.600 85.800 141.000 86.200 ;
        RECT 157.400 85.800 157.800 86.200 ;
        RECT 165.400 86.100 165.800 86.200 ;
        RECT 165.400 85.800 166.500 86.100 ;
        RECT 7.800 85.200 8.100 85.800 ;
        RECT 104.600 85.200 104.900 85.800 ;
        RECT 7.800 84.800 8.200 85.200 ;
        RECT 35.800 85.100 36.200 85.200 ;
        RECT 37.400 85.100 37.800 85.200 ;
        RECT 35.800 84.800 41.700 85.100 ;
        RECT 41.400 84.200 41.700 84.800 ;
        RECT 43.000 84.800 43.400 85.200 ;
        RECT 46.200 85.100 46.600 85.200 ;
        RECT 47.800 85.100 48.200 85.200 ;
        RECT 46.200 84.800 48.200 85.100 ;
        RECT 104.600 84.800 105.000 85.200 ;
        RECT 138.200 85.100 138.600 85.200 ;
        RECT 140.600 85.100 140.900 85.800 ;
        RECT 138.200 84.800 140.900 85.100 ;
        RECT 166.200 85.200 166.500 85.800 ;
        RECT 166.200 84.800 166.600 85.200 ;
        RECT 167.800 85.100 168.200 85.200 ;
        RECT 175.000 85.100 175.400 85.200 ;
        RECT 183.800 85.100 184.200 85.200 ;
        RECT 167.800 84.800 184.200 85.100 ;
        RECT 41.400 83.800 41.800 84.200 ;
        RECT 43.000 84.100 43.300 84.800 ;
        RECT 59.000 84.100 59.400 84.200 ;
        RECT 43.000 83.800 59.400 84.100 ;
        RECT 137.400 84.100 137.800 84.200 ;
        RECT 139.800 84.100 140.200 84.200 ;
        RECT 137.400 83.800 140.200 84.100 ;
        RECT 168.600 84.100 169.000 84.200 ;
        RECT 171.000 84.100 171.400 84.200 ;
        RECT 168.600 83.800 171.400 84.100 ;
        RECT 25.400 83.100 25.800 83.200 ;
        RECT 86.200 83.100 86.600 83.200 ;
        RECT 25.400 82.800 86.600 83.100 ;
        RECT 164.600 83.100 165.000 83.200 ;
        RECT 173.400 83.100 173.800 83.200 ;
        RECT 178.200 83.100 178.600 83.200 ;
        RECT 186.200 83.100 186.600 83.200 ;
        RECT 164.600 82.800 186.600 83.100 ;
        RECT 15.000 82.100 15.400 82.200 ;
        RECT 16.600 82.100 17.000 82.200 ;
        RECT 15.000 81.800 17.000 82.100 ;
        RECT 28.600 82.100 29.000 82.200 ;
        RECT 33.400 82.100 33.800 82.200 ;
        RECT 50.200 82.100 50.600 82.200 ;
        RECT 28.600 81.800 50.600 82.100 ;
        RECT 71.800 82.100 72.200 82.200 ;
        RECT 80.600 82.100 81.000 82.200 ;
        RECT 100.600 82.100 101.000 82.200 ;
        RECT 119.800 82.100 120.200 82.200 ;
        RECT 71.800 81.800 120.200 82.100 ;
        RECT 162.200 82.100 162.600 82.200 ;
        RECT 165.400 82.100 165.800 82.200 ;
        RECT 171.000 82.100 171.400 82.200 ;
        RECT 162.200 81.800 171.400 82.100 ;
        RECT 34.200 81.100 34.600 81.200 ;
        RECT 42.200 81.100 42.600 81.200 ;
        RECT 34.200 80.800 42.600 81.100 ;
        RECT 98.200 81.100 98.600 81.200 ;
        RECT 107.800 81.100 108.200 81.200 ;
        RECT 98.200 80.800 108.200 81.100 ;
        RECT 10.200 80.100 10.600 80.200 ;
        RECT 11.800 80.100 12.200 80.200 ;
        RECT 10.200 79.800 12.200 80.100 ;
        RECT 86.200 80.100 86.600 80.200 ;
        RECT 88.600 80.100 89.000 80.200 ;
        RECT 99.000 80.100 99.400 80.200 ;
        RECT 86.200 79.800 99.400 80.100 ;
        RECT 6.200 79.100 6.600 79.200 ;
        RECT 9.400 79.100 9.800 79.200 ;
        RECT 6.200 78.800 9.800 79.100 ;
        RECT 38.200 79.100 38.600 79.200 ;
        RECT 39.000 79.100 39.400 79.200 ;
        RECT 38.200 78.800 39.400 79.100 ;
        RECT 39.800 79.100 40.200 79.200 ;
        RECT 99.800 79.100 100.200 79.200 ;
        RECT 114.200 79.100 114.600 79.200 ;
        RECT 39.800 78.800 114.600 79.100 ;
        RECT 117.400 79.100 117.800 79.200 ;
        RECT 121.400 79.100 121.800 79.200 ;
        RECT 117.400 78.800 121.800 79.100 ;
        RECT 83.000 78.100 83.400 78.200 ;
        RECT 86.200 78.100 86.600 78.200 ;
        RECT 89.400 78.100 89.800 78.200 ;
        RECT 137.400 78.100 137.800 78.200 ;
        RECT 83.000 77.800 137.800 78.100 ;
        RECT 31.800 77.100 32.200 77.200 ;
        RECT 45.400 77.100 45.800 77.200 ;
        RECT 48.600 77.100 49.000 77.200 ;
        RECT 31.800 76.800 49.000 77.100 ;
        RECT 55.800 76.800 56.200 77.200 ;
        RECT 65.400 77.100 65.800 77.200 ;
        RECT 78.200 77.100 78.600 77.200 ;
        RECT 65.400 76.800 78.600 77.100 ;
        RECT 166.200 77.100 166.600 77.200 ;
        RECT 173.400 77.100 173.800 77.200 ;
        RECT 166.200 76.800 173.800 77.100 ;
        RECT 178.200 77.100 178.600 77.200 ;
        RECT 180.600 77.100 181.000 77.200 ;
        RECT 178.200 76.800 181.000 77.100 ;
        RECT 31.000 76.100 31.400 76.200 ;
        RECT 40.600 76.100 41.000 76.200 ;
        RECT 31.000 75.800 41.000 76.100 ;
        RECT 43.000 76.100 43.400 76.200 ;
        RECT 51.000 76.100 51.400 76.200 ;
        RECT 53.400 76.100 53.800 76.200 ;
        RECT 43.000 75.800 53.800 76.100 ;
        RECT 55.800 76.100 56.100 76.800 ;
        RECT 65.400 76.100 65.800 76.200 ;
        RECT 55.800 75.800 65.800 76.100 ;
        RECT 77.400 75.800 77.800 76.200 ;
        RECT 78.200 76.100 78.600 76.200 ;
        RECT 81.400 76.100 81.800 76.200 ;
        RECT 78.200 75.800 81.800 76.100 ;
        RECT 83.800 76.100 84.200 76.200 ;
        RECT 88.600 76.100 89.000 76.200 ;
        RECT 83.800 75.800 89.000 76.100 ;
        RECT 91.800 76.100 92.200 76.200 ;
        RECT 103.000 76.100 103.400 76.200 ;
        RECT 91.800 75.800 103.400 76.100 ;
        RECT 121.400 76.100 121.800 76.200 ;
        RECT 127.000 76.100 127.400 76.200 ;
        RECT 121.400 75.800 127.400 76.100 ;
        RECT 164.600 76.100 165.000 76.200 ;
        RECT 166.200 76.100 166.600 76.200 ;
        RECT 164.600 75.800 166.600 76.100 ;
        RECT 168.600 76.100 169.000 76.200 ;
        RECT 170.200 76.100 170.600 76.200 ;
        RECT 168.600 75.800 170.600 76.100 ;
        RECT 179.800 75.800 180.200 76.200 ;
        RECT 77.400 75.200 77.700 75.800 ;
        RECT 5.400 75.100 5.800 75.200 ;
        RECT 7.000 75.100 7.400 75.200 ;
        RECT 5.400 74.800 7.400 75.100 ;
        RECT 9.400 75.100 9.800 75.200 ;
        RECT 16.600 75.100 17.000 75.200 ;
        RECT 42.200 75.100 42.600 75.200 ;
        RECT 9.400 74.800 17.000 75.100 ;
        RECT 37.400 74.800 42.600 75.100 ;
        RECT 47.800 75.100 48.200 75.200 ;
        RECT 56.600 75.100 57.000 75.200 ;
        RECT 47.800 74.800 57.000 75.100 ;
        RECT 59.800 75.100 60.200 75.200 ;
        RECT 76.600 75.100 77.000 75.200 ;
        RECT 59.800 74.800 77.000 75.100 ;
        RECT 77.400 74.800 77.800 75.200 ;
        RECT 79.800 75.100 80.200 75.200 ;
        RECT 81.400 75.100 81.800 75.200 ;
        RECT 79.800 74.800 81.800 75.100 ;
        RECT 84.600 75.100 85.000 75.200 ;
        RECT 85.400 75.100 85.800 75.200 ;
        RECT 84.600 74.800 85.800 75.100 ;
        RECT 87.800 75.100 88.200 75.200 ;
        RECT 92.600 75.100 93.000 75.200 ;
        RECT 98.200 75.100 98.600 75.200 ;
        RECT 87.800 74.800 98.600 75.100 ;
        RECT 125.400 75.100 125.800 75.200 ;
        RECT 126.200 75.100 126.600 75.200 ;
        RECT 125.400 74.800 126.600 75.100 ;
        RECT 159.000 75.100 159.400 75.200 ;
        RECT 164.600 75.100 165.000 75.200 ;
        RECT 166.200 75.100 166.600 75.200 ;
        RECT 159.000 74.800 166.600 75.100 ;
        RECT 174.200 75.100 174.600 75.200 ;
        RECT 179.800 75.100 180.100 75.800 ;
        RECT 174.200 74.800 180.100 75.100 ;
        RECT 185.400 74.800 185.800 75.200 ;
        RECT 37.400 74.700 37.800 74.800 ;
        RECT 7.000 74.100 7.400 74.200 ;
        RECT 14.200 74.100 14.600 74.200 ;
        RECT 7.000 73.800 14.600 74.100 ;
        RECT 36.600 74.100 37.000 74.200 ;
        RECT 39.800 74.100 40.200 74.200 ;
        RECT 43.000 74.100 43.400 74.200 ;
        RECT 55.800 74.100 56.200 74.200 ;
        RECT 57.400 74.100 57.800 74.200 ;
        RECT 36.600 73.800 43.400 74.100 ;
        RECT 50.200 73.800 57.800 74.100 ;
        RECT 63.000 73.800 63.400 74.200 ;
        RECT 76.600 74.100 77.000 74.200 ;
        RECT 80.600 74.100 81.000 74.200 ;
        RECT 86.200 74.100 86.600 74.200 ;
        RECT 88.600 74.100 89.000 74.200 ;
        RECT 76.600 73.800 89.000 74.100 ;
        RECT 111.000 74.100 111.400 74.200 ;
        RECT 116.600 74.100 117.000 74.200 ;
        RECT 111.000 73.800 117.000 74.100 ;
        RECT 134.200 74.100 134.600 74.200 ;
        RECT 136.600 74.100 137.000 74.200 ;
        RECT 137.400 74.100 137.800 74.200 ;
        RECT 134.200 73.800 137.800 74.100 ;
        RECT 146.200 74.100 146.600 74.200 ;
        RECT 146.200 73.800 155.300 74.100 ;
        RECT 50.200 73.200 50.500 73.800 ;
        RECT 9.400 73.100 9.800 73.200 ;
        RECT 28.600 73.100 29.000 73.200 ;
        RECT 39.800 73.100 40.200 73.200 ;
        RECT 9.400 72.800 40.200 73.100 ;
        RECT 47.800 73.100 48.200 73.200 ;
        RECT 50.200 73.100 50.600 73.200 ;
        RECT 47.800 72.800 50.600 73.100 ;
        RECT 51.800 73.100 52.200 73.200 ;
        RECT 53.400 73.100 53.800 73.200 ;
        RECT 51.800 72.800 53.800 73.100 ;
        RECT 57.400 73.100 57.800 73.200 ;
        RECT 59.800 73.100 60.200 73.200 ;
        RECT 57.400 72.800 60.200 73.100 ;
        RECT 63.000 73.100 63.300 73.800 ;
        RECT 63.800 73.100 64.200 73.200 ;
        RECT 63.000 72.800 64.200 73.100 ;
        RECT 73.400 73.100 73.800 73.200 ;
        RECT 79.800 73.100 80.200 73.200 ;
        RECT 107.000 73.100 107.400 73.200 ;
        RECT 109.400 73.100 109.800 73.200 ;
        RECT 125.400 73.100 125.800 73.200 ;
        RECT 73.400 72.800 78.500 73.100 ;
        RECT 79.800 72.800 83.300 73.100 ;
        RECT 107.000 72.800 125.800 73.100 ;
        RECT 127.800 73.100 128.200 73.200 ;
        RECT 134.200 73.100 134.500 73.800 ;
        RECT 155.000 73.200 155.300 73.800 ;
        RECT 163.000 73.800 163.400 74.200 ;
        RECT 164.600 74.100 165.000 74.200 ;
        RECT 167.000 74.100 167.400 74.200 ;
        RECT 164.600 73.800 167.400 74.100 ;
        RECT 184.600 74.100 185.000 74.200 ;
        RECT 185.400 74.100 185.700 74.800 ;
        RECT 184.600 73.800 185.700 74.100 ;
        RECT 127.800 72.800 134.500 73.100 ;
        RECT 151.800 73.100 152.200 73.200 ;
        RECT 151.800 72.800 152.900 73.100 ;
        RECT 155.000 72.800 155.400 73.200 ;
        RECT 163.000 73.100 163.300 73.800 ;
        RECT 169.400 73.100 169.800 73.200 ;
        RECT 163.000 72.800 169.800 73.100 ;
        RECT 171.000 73.100 171.400 73.200 ;
        RECT 175.800 73.100 176.200 73.200 ;
        RECT 171.000 72.800 176.200 73.100 ;
        RECT 78.200 72.200 78.500 72.800 ;
        RECT 83.000 72.200 83.300 72.800 ;
        RECT 152.600 72.200 152.900 72.800 ;
        RECT 23.000 72.100 23.400 72.200 ;
        RECT 30.200 72.100 30.600 72.200 ;
        RECT 23.000 71.800 30.600 72.100 ;
        RECT 64.600 72.100 65.000 72.200 ;
        RECT 70.200 72.100 70.600 72.200 ;
        RECT 64.600 71.800 70.600 72.100 ;
        RECT 78.200 71.800 78.600 72.200 ;
        RECT 83.000 71.800 83.400 72.200 ;
        RECT 96.600 72.100 97.000 72.200 ;
        RECT 108.600 72.100 109.000 72.200 ;
        RECT 111.000 72.100 111.400 72.200 ;
        RECT 96.600 71.800 111.400 72.100 ;
        RECT 152.600 71.800 153.000 72.200 ;
        RECT 165.400 72.100 165.800 72.200 ;
        RECT 167.800 72.100 168.200 72.200 ;
        RECT 165.400 71.800 168.200 72.100 ;
        RECT 42.200 71.100 42.600 71.200 ;
        RECT 62.200 71.100 62.600 71.200 ;
        RECT 42.200 70.800 62.600 71.100 ;
        RECT 63.000 71.100 63.400 71.200 ;
        RECT 86.200 71.100 86.600 71.200 ;
        RECT 63.000 70.800 86.600 71.100 ;
        RECT 163.800 71.100 164.200 71.200 ;
        RECT 177.400 71.100 177.800 71.200 ;
        RECT 163.800 70.800 177.800 71.100 ;
        RECT 38.200 70.100 38.600 70.200 ;
        RECT 53.400 70.100 53.800 70.200 ;
        RECT 63.000 70.100 63.400 70.200 ;
        RECT 67.000 70.100 67.400 70.200 ;
        RECT 38.200 69.800 67.400 70.100 ;
        RECT 77.400 70.100 77.800 70.200 ;
        RECT 95.800 70.100 96.200 70.200 ;
        RECT 77.400 69.800 96.200 70.100 ;
        RECT 139.800 70.100 140.200 70.200 ;
        RECT 147.800 70.100 148.200 70.200 ;
        RECT 139.800 69.800 148.200 70.100 ;
        RECT 173.400 70.100 173.800 70.200 ;
        RECT 192.600 70.100 193.000 70.200 ;
        RECT 173.400 69.800 193.000 70.100 ;
        RECT 77.400 69.200 77.700 69.800 ;
        RECT 62.200 69.100 62.600 69.200 ;
        RECT 63.000 69.100 63.400 69.200 ;
        RECT 62.200 68.800 63.400 69.100 ;
        RECT 77.400 68.800 77.800 69.200 ;
        RECT 79.000 69.100 79.400 69.200 ;
        RECT 87.800 69.100 88.200 69.200 ;
        RECT 79.000 68.800 88.200 69.100 ;
        RECT 88.600 69.100 89.000 69.200 ;
        RECT 94.200 69.100 94.600 69.200 ;
        RECT 88.600 68.800 94.600 69.100 ;
        RECT 95.800 69.100 96.100 69.800 ;
        RECT 97.400 69.100 97.800 69.200 ;
        RECT 95.800 68.800 97.800 69.100 ;
        RECT 116.600 69.100 117.000 69.200 ;
        RECT 133.400 69.100 133.800 69.200 ;
        RECT 116.600 68.800 133.800 69.100 ;
        RECT 155.000 69.100 155.400 69.200 ;
        RECT 166.200 69.100 166.600 69.200 ;
        RECT 155.000 68.800 166.600 69.100 ;
        RECT 179.000 68.800 179.400 69.200 ;
        RECT 183.800 69.100 184.200 69.200 ;
        RECT 187.800 69.100 188.200 69.200 ;
        RECT 193.400 69.100 193.800 69.200 ;
        RECT 183.800 68.800 193.800 69.100 ;
        RECT 52.600 68.100 53.000 68.200 ;
        RECT 55.000 68.100 55.400 68.200 ;
        RECT 63.800 68.100 64.200 68.200 ;
        RECT 52.600 67.800 64.200 68.100 ;
        RECT 71.000 68.100 71.400 68.200 ;
        RECT 82.200 68.100 82.600 68.200 ;
        RECT 87.800 68.100 88.200 68.200 ;
        RECT 93.400 68.100 93.800 68.200 ;
        RECT 71.000 67.800 93.800 68.100 ;
        RECT 113.400 68.100 113.800 68.200 ;
        RECT 123.800 68.100 124.200 68.200 ;
        RECT 160.600 68.100 161.000 68.200 ;
        RECT 113.400 67.800 161.000 68.100 ;
        RECT 169.400 68.100 169.800 68.200 ;
        RECT 179.000 68.100 179.300 68.800 ;
        RECT 169.400 67.800 179.300 68.100 ;
        RECT 180.600 67.800 181.000 68.200 ;
        RECT 27.000 67.100 27.400 67.200 ;
        RECT 37.400 67.100 37.800 67.200 ;
        RECT 18.200 66.800 37.800 67.100 ;
        RECT 54.200 66.800 54.600 67.200 ;
        RECT 69.400 67.100 69.800 67.200 ;
        RECT 73.400 67.100 73.800 67.200 ;
        RECT 69.400 66.800 73.800 67.100 ;
        RECT 76.600 67.100 77.000 67.200 ;
        RECT 79.800 67.100 80.200 67.200 ;
        RECT 76.600 66.800 80.200 67.100 ;
        RECT 91.800 66.800 92.200 67.200 ;
        RECT 94.200 67.100 94.600 67.200 ;
        RECT 103.800 67.100 104.200 67.200 ;
        RECT 94.200 66.800 104.200 67.100 ;
        RECT 107.000 66.800 107.400 67.200 ;
        RECT 155.000 67.100 155.400 67.200 ;
        RECT 159.000 67.100 159.400 67.200 ;
        RECT 155.000 66.800 159.400 67.100 ;
        RECT 163.000 67.100 163.400 67.200 ;
        RECT 164.600 67.100 165.000 67.200 ;
        RECT 163.000 66.800 165.000 67.100 ;
        RECT 166.200 67.100 166.600 67.200 ;
        RECT 180.600 67.100 180.900 67.800 ;
        RECT 166.200 66.800 180.900 67.100 ;
        RECT 182.200 67.100 182.600 67.200 ;
        RECT 187.000 67.100 187.400 67.200 ;
        RECT 182.200 66.800 187.400 67.100 ;
        RECT 18.200 66.200 18.500 66.800 ;
        RECT 18.200 65.800 18.600 66.200 ;
        RECT 41.400 66.100 41.800 66.200 ;
        RECT 43.000 66.100 43.400 66.200 ;
        RECT 50.200 66.100 50.600 66.200 ;
        RECT 54.200 66.100 54.500 66.800 ;
        RECT 41.400 65.800 54.500 66.100 ;
        RECT 56.600 66.100 57.000 66.200 ;
        RECT 59.800 66.100 60.200 66.200 ;
        RECT 56.600 65.800 60.200 66.100 ;
        RECT 83.000 66.100 83.400 66.300 ;
        RECT 87.800 66.100 88.200 66.200 ;
        RECT 91.800 66.100 92.100 66.800 ;
        RECT 83.000 65.800 92.100 66.100 ;
        RECT 107.000 66.200 107.300 66.800 ;
        RECT 159.000 66.200 159.300 66.800 ;
        RECT 107.000 65.800 107.400 66.200 ;
        RECT 135.000 66.100 135.400 66.200 ;
        RECT 142.200 66.100 142.600 66.200 ;
        RECT 147.000 66.100 147.400 66.200 ;
        RECT 154.200 66.100 154.600 66.200 ;
        RECT 135.000 65.800 147.400 66.100 ;
        RECT 153.400 65.800 154.600 66.100 ;
        RECT 159.000 65.800 159.400 66.200 ;
        RECT 170.200 66.100 170.600 66.200 ;
        RECT 171.000 66.100 171.400 66.200 ;
        RECT 170.200 65.800 171.400 66.100 ;
        RECT 174.200 66.100 174.600 66.200 ;
        RECT 175.000 66.100 175.400 66.200 ;
        RECT 174.200 65.800 175.400 66.100 ;
        RECT 178.200 66.100 178.600 66.200 ;
        RECT 182.200 66.100 182.500 66.800 ;
        RECT 178.200 65.800 182.500 66.100 ;
        RECT 15.800 65.100 16.200 65.200 ;
        RECT 28.600 65.100 29.000 65.200 ;
        RECT 33.400 65.100 33.800 65.200 ;
        RECT 15.800 64.800 20.100 65.100 ;
        RECT 28.600 64.800 33.800 65.100 ;
        RECT 47.800 65.100 48.200 65.200 ;
        RECT 53.400 65.100 53.800 65.200 ;
        RECT 59.000 65.100 59.400 65.200 ;
        RECT 47.800 64.800 59.400 65.100 ;
        RECT 164.600 65.100 165.000 65.200 ;
        RECT 173.400 65.100 173.800 65.200 ;
        RECT 164.600 64.800 173.800 65.100 ;
        RECT 19.800 64.200 20.100 64.800 ;
        RECT 19.800 63.800 20.200 64.200 ;
        RECT 27.800 64.100 28.200 64.200 ;
        RECT 84.600 64.100 85.000 64.200 ;
        RECT 122.200 64.100 122.600 64.200 ;
        RECT 124.600 64.100 125.000 64.200 ;
        RECT 27.800 63.800 125.000 64.100 ;
        RECT 159.800 64.100 160.200 64.200 ;
        RECT 163.000 64.100 163.400 64.200 ;
        RECT 169.400 64.100 169.800 64.200 ;
        RECT 159.800 63.800 169.800 64.100 ;
        RECT 160.600 63.100 161.000 63.200 ;
        RECT 162.200 63.100 162.600 63.200 ;
        RECT 171.800 63.100 172.200 63.200 ;
        RECT 160.600 62.800 172.200 63.100 ;
        RECT 18.200 62.100 18.600 62.200 ;
        RECT 22.200 62.100 22.600 62.200 ;
        RECT 29.400 62.100 29.800 62.200 ;
        RECT 36.600 62.100 37.000 62.200 ;
        RECT 18.200 61.800 37.000 62.100 ;
        RECT 35.000 60.100 35.400 60.200 ;
        RECT 38.200 60.100 38.600 60.200 ;
        RECT 35.000 59.800 38.600 60.100 ;
        RECT 193.400 59.800 193.800 60.200 ;
        RECT 193.400 59.200 193.700 59.800 ;
        RECT 69.400 59.100 69.800 59.200 ;
        RECT 73.400 59.100 73.800 59.200 ;
        RECT 69.400 58.800 73.800 59.100 ;
        RECT 193.400 58.800 193.800 59.200 ;
        RECT 51.000 58.100 51.400 58.200 ;
        RECT 80.600 58.100 81.000 58.200 ;
        RECT 51.000 57.800 81.000 58.100 ;
        RECT 139.800 58.100 140.200 58.200 ;
        RECT 140.600 58.100 141.000 58.200 ;
        RECT 149.400 58.100 149.800 58.200 ;
        RECT 163.800 58.100 164.200 58.200 ;
        RECT 139.800 57.800 164.200 58.100 ;
        RECT 167.000 58.100 167.400 58.200 ;
        RECT 169.400 58.100 169.800 58.200 ;
        RECT 170.200 58.100 170.600 58.200 ;
        RECT 167.000 57.800 170.600 58.100 ;
        RECT 9.400 57.100 9.800 57.200 ;
        RECT 19.800 57.100 20.200 57.200 ;
        RECT 25.400 57.100 25.800 57.200 ;
        RECT 9.400 56.800 12.900 57.100 ;
        RECT 19.800 56.800 25.800 57.100 ;
        RECT 47.800 57.100 48.200 57.200 ;
        RECT 72.600 57.100 73.000 57.200 ;
        RECT 75.800 57.100 76.200 57.200 ;
        RECT 47.800 56.800 76.200 57.100 ;
        RECT 80.600 56.800 81.000 57.200 ;
        RECT 105.400 57.100 105.800 57.200 ;
        RECT 110.200 57.100 110.600 57.200 ;
        RECT 105.400 56.800 110.600 57.100 ;
        RECT 115.800 56.800 116.200 57.200 ;
        RECT 147.800 57.100 148.200 57.200 ;
        RECT 178.200 57.100 178.600 57.200 ;
        RECT 185.400 57.100 185.800 57.200 ;
        RECT 186.200 57.100 186.600 57.200 ;
        RECT 147.800 56.800 169.700 57.100 ;
        RECT 178.200 56.800 186.600 57.100 ;
        RECT 12.600 56.200 12.900 56.800 ;
        RECT 80.600 56.200 80.900 56.800 ;
        RECT 8.600 56.100 9.000 56.200 ;
        RECT 10.200 56.100 10.600 56.200 ;
        RECT 8.600 55.800 10.600 56.100 ;
        RECT 12.600 55.800 13.000 56.200 ;
        RECT 23.000 55.800 23.400 56.200 ;
        RECT 31.800 56.100 32.200 56.200 ;
        RECT 35.800 56.100 36.200 56.200 ;
        RECT 31.800 55.800 36.200 56.100 ;
        RECT 37.400 56.100 37.800 56.200 ;
        RECT 39.800 56.100 40.200 56.200 ;
        RECT 44.600 56.100 45.000 56.200 ;
        RECT 37.400 55.800 45.000 56.100 ;
        RECT 45.400 56.100 45.800 56.200 ;
        RECT 49.400 56.100 49.800 56.200 ;
        RECT 51.800 56.100 52.200 56.200 ;
        RECT 61.400 56.100 61.800 56.200 ;
        RECT 76.600 56.100 77.000 56.200 ;
        RECT 45.400 55.800 77.000 56.100 ;
        RECT 80.600 55.800 81.000 56.200 ;
        RECT 83.800 56.100 84.200 56.200 ;
        RECT 86.200 56.100 86.600 56.200 ;
        RECT 83.000 55.800 86.600 56.100 ;
        RECT 87.000 56.100 87.400 56.200 ;
        RECT 103.800 56.100 104.200 56.200 ;
        RECT 87.000 55.800 104.200 56.100 ;
        RECT 105.400 56.100 105.800 56.200 ;
        RECT 111.800 56.100 112.200 56.200 ;
        RECT 115.800 56.100 116.100 56.800 ;
        RECT 169.400 56.200 169.700 56.800 ;
        RECT 163.000 56.100 163.400 56.200 ;
        RECT 105.400 55.800 116.100 56.100 ;
        RECT 160.600 55.800 163.400 56.100 ;
        RECT 169.400 56.100 169.800 56.200 ;
        RECT 171.000 56.100 171.400 56.200 ;
        RECT 169.400 55.800 171.400 56.100 ;
        RECT 171.800 56.100 172.200 56.200 ;
        RECT 179.800 56.100 180.200 56.200 ;
        RECT 171.800 55.800 180.200 56.100 ;
        RECT 10.200 55.100 10.500 55.800 ;
        RECT 23.000 55.100 23.300 55.800 ;
        RECT 160.600 55.200 160.900 55.800 ;
        RECT 47.800 55.100 48.200 55.200 ;
        RECT 10.200 54.800 48.200 55.100 ;
        RECT 48.600 55.100 49.000 55.200 ;
        RECT 51.000 55.100 51.400 55.200 ;
        RECT 71.000 55.100 71.400 55.200 ;
        RECT 48.600 54.800 51.400 55.100 ;
        RECT 57.400 54.800 71.400 55.100 ;
        RECT 75.800 55.100 76.200 55.200 ;
        RECT 87.800 55.100 88.200 55.200 ;
        RECT 75.800 54.800 88.200 55.100 ;
        RECT 108.600 55.100 109.000 55.200 ;
        RECT 112.600 55.100 113.000 55.200 ;
        RECT 114.200 55.100 114.600 55.200 ;
        RECT 108.600 54.800 113.000 55.100 ;
        RECT 113.400 54.800 114.600 55.100 ;
        RECT 117.400 55.100 117.800 55.200 ;
        RECT 121.400 55.100 121.800 55.200 ;
        RECT 117.400 54.800 121.800 55.100 ;
        RECT 145.400 55.100 145.800 55.200 ;
        RECT 147.000 55.100 147.400 55.200 ;
        RECT 145.400 54.800 147.400 55.100 ;
        RECT 152.600 55.100 153.000 55.200 ;
        RECT 152.600 54.800 159.300 55.100 ;
        RECT 160.600 54.800 161.000 55.200 ;
        RECT 167.000 55.100 167.400 55.200 ;
        RECT 175.800 55.100 176.200 55.200 ;
        RECT 167.000 54.800 176.200 55.100 ;
        RECT 177.400 55.100 177.800 55.200 ;
        RECT 179.800 55.100 180.200 55.200 ;
        RECT 177.400 54.800 180.200 55.100 ;
        RECT 57.400 54.700 57.800 54.800 ;
        RECT 67.000 54.700 67.400 54.800 ;
        RECT 159.000 54.200 159.300 54.800 ;
        RECT 11.000 54.100 11.400 54.200 ;
        RECT 14.200 54.100 14.600 54.200 ;
        RECT 11.000 53.800 14.600 54.100 ;
        RECT 22.200 54.100 22.600 54.200 ;
        RECT 24.600 54.100 25.000 54.200 ;
        RECT 22.200 53.800 25.000 54.100 ;
        RECT 58.200 54.100 58.600 54.200 ;
        RECT 64.600 54.100 65.000 54.200 ;
        RECT 58.200 53.800 65.000 54.100 ;
        RECT 72.600 54.100 73.000 54.200 ;
        RECT 77.400 54.100 77.800 54.200 ;
        RECT 72.600 53.800 77.800 54.100 ;
        RECT 83.800 54.100 84.200 54.200 ;
        RECT 84.600 54.100 85.000 54.200 ;
        RECT 83.800 53.800 85.000 54.100 ;
        RECT 87.800 54.100 88.200 54.200 ;
        RECT 108.600 54.100 109.000 54.200 ;
        RECT 109.400 54.100 109.800 54.200 ;
        RECT 118.200 54.100 118.600 54.200 ;
        RECT 87.800 53.800 118.600 54.100 ;
        RECT 119.000 54.100 119.400 54.200 ;
        RECT 119.800 54.100 120.200 54.200 ;
        RECT 119.000 53.800 120.200 54.100 ;
        RECT 120.600 54.100 121.000 54.200 ;
        RECT 130.200 54.100 130.600 54.200 ;
        RECT 120.600 53.800 130.600 54.100 ;
        RECT 159.000 53.800 159.400 54.200 ;
        RECT 167.800 54.100 168.200 54.200 ;
        RECT 171.000 54.100 171.400 54.200 ;
        RECT 167.800 53.800 171.400 54.100 ;
        RECT 172.600 54.100 173.000 54.200 ;
        RECT 176.600 54.100 177.000 54.200 ;
        RECT 178.200 54.100 178.600 54.200 ;
        RECT 172.600 53.800 178.600 54.100 ;
        RECT 179.000 54.100 179.400 54.200 ;
        RECT 182.200 54.100 182.600 54.200 ;
        RECT 179.000 53.800 182.600 54.100 ;
        RECT 23.800 53.100 24.200 53.200 ;
        RECT 27.800 53.100 28.200 53.200 ;
        RECT 30.200 53.100 30.600 53.200 ;
        RECT 23.800 52.800 30.600 53.100 ;
        RECT 42.200 53.100 42.600 53.200 ;
        RECT 47.800 53.100 48.200 53.200 ;
        RECT 42.200 52.800 48.200 53.100 ;
        RECT 57.400 53.100 57.800 53.200 ;
        RECT 72.600 53.100 73.000 53.200 ;
        RECT 83.800 53.100 84.200 53.200 ;
        RECT 57.400 52.800 84.200 53.100 ;
        RECT 86.200 53.100 86.600 53.200 ;
        RECT 87.000 53.100 87.400 53.200 ;
        RECT 86.200 52.800 87.400 53.100 ;
        RECT 90.200 53.100 90.600 53.200 ;
        RECT 93.400 53.100 93.800 53.200 ;
        RECT 90.200 52.800 93.800 53.100 ;
        RECT 103.000 53.100 103.400 53.200 ;
        RECT 113.400 53.100 113.800 53.200 ;
        RECT 103.000 52.800 113.800 53.100 ;
        RECT 115.000 53.100 115.400 53.200 ;
        RECT 136.600 53.100 137.000 53.200 ;
        RECT 115.000 52.800 137.000 53.100 ;
        RECT 151.800 53.100 152.200 53.200 ;
        RECT 155.800 53.100 156.200 53.200 ;
        RECT 151.800 52.800 156.200 53.100 ;
        RECT 161.400 53.100 161.800 53.200 ;
        RECT 172.600 53.100 173.000 53.200 ;
        RECT 161.400 52.800 173.000 53.100 ;
        RECT 193.400 53.100 193.800 53.200 ;
        RECT 194.200 53.100 194.600 53.200 ;
        RECT 193.400 52.800 194.600 53.100 ;
        RECT 71.000 52.200 71.300 52.800 ;
        RECT 71.000 51.800 71.400 52.200 ;
        RECT 83.800 52.100 84.200 52.200 ;
        RECT 98.200 52.100 98.600 52.200 ;
        RECT 83.800 51.800 98.600 52.100 ;
        RECT 114.200 52.100 114.600 52.200 ;
        RECT 123.800 52.100 124.200 52.200 ;
        RECT 114.200 51.800 124.200 52.100 ;
        RECT 156.600 52.100 157.000 52.200 ;
        RECT 165.400 52.100 165.800 52.200 ;
        RECT 156.600 51.800 165.800 52.100 ;
        RECT 111.800 51.100 112.200 51.200 ;
        RECT 139.000 51.100 139.400 51.200 ;
        RECT 159.800 51.100 160.200 51.200 ;
        RECT 111.800 50.800 160.200 51.100 ;
        RECT 18.200 50.100 18.600 50.200 ;
        RECT 21.400 50.100 21.800 50.200 ;
        RECT 27.800 50.100 28.200 50.200 ;
        RECT 18.200 49.800 28.200 50.100 ;
        RECT 33.400 49.800 33.800 50.200 ;
        RECT 38.200 49.800 38.600 50.200 ;
        RECT 40.600 50.100 41.000 50.200 ;
        RECT 43.000 50.100 43.400 50.200 ;
        RECT 40.600 49.800 43.400 50.100 ;
        RECT 79.000 49.800 79.400 50.200 ;
        RECT 88.600 49.800 89.000 50.200 ;
        RECT 162.200 50.100 162.600 50.200 ;
        RECT 168.600 50.100 169.000 50.200 ;
        RECT 162.200 49.800 169.000 50.100 ;
        RECT 171.800 50.100 172.200 50.200 ;
        RECT 180.600 50.100 181.000 50.200 ;
        RECT 171.800 49.800 181.000 50.100 ;
        RECT 3.800 49.100 4.200 49.200 ;
        RECT 11.000 49.100 11.400 49.200 ;
        RECT 28.600 49.100 29.000 49.200 ;
        RECT 3.800 48.800 29.000 49.100 ;
        RECT 30.200 49.100 30.600 49.200 ;
        RECT 33.400 49.100 33.700 49.800 ;
        RECT 30.200 48.800 33.700 49.100 ;
        RECT 38.200 49.200 38.500 49.800 ;
        RECT 79.000 49.200 79.300 49.800 ;
        RECT 88.600 49.200 88.900 49.800 ;
        RECT 38.200 48.800 38.600 49.200 ;
        RECT 39.000 49.100 39.400 49.200 ;
        RECT 43.000 49.100 43.400 49.200 ;
        RECT 39.000 48.800 43.400 49.100 ;
        RECT 48.600 49.100 49.000 49.200 ;
        RECT 68.600 49.100 69.000 49.200 ;
        RECT 48.600 48.800 69.000 49.100 ;
        RECT 79.000 48.800 79.400 49.200 ;
        RECT 88.600 48.800 89.000 49.200 ;
        RECT 100.600 49.100 101.000 49.200 ;
        RECT 119.000 49.100 119.400 49.200 ;
        RECT 137.400 49.100 137.800 49.200 ;
        RECT 99.800 48.800 137.800 49.100 ;
        RECT 139.800 49.100 140.200 49.200 ;
        RECT 152.600 49.100 153.000 49.200 ;
        RECT 139.800 48.800 153.000 49.100 ;
        RECT 159.000 49.100 159.400 49.200 ;
        RECT 164.600 49.100 165.000 49.200 ;
        RECT 180.600 49.100 181.000 49.200 ;
        RECT 183.800 49.100 184.200 49.200 ;
        RECT 159.000 48.800 184.200 49.100 ;
        RECT 8.600 48.100 9.000 48.200 ;
        RECT 13.400 48.100 13.800 48.200 ;
        RECT 15.800 48.100 16.200 48.200 ;
        RECT 8.600 47.800 16.200 48.100 ;
        RECT 30.200 48.100 30.600 48.200 ;
        RECT 55.800 48.100 56.200 48.200 ;
        RECT 30.200 47.800 56.200 48.100 ;
        RECT 67.800 48.100 68.200 48.200 ;
        RECT 68.600 48.100 69.000 48.200 ;
        RECT 67.800 47.800 69.000 48.100 ;
        RECT 80.600 48.100 81.000 48.200 ;
        RECT 83.000 48.100 83.400 48.200 ;
        RECT 90.200 48.100 90.600 48.200 ;
        RECT 106.200 48.100 106.600 48.200 ;
        RECT 80.600 47.800 106.600 48.100 ;
        RECT 143.800 48.100 144.200 48.200 ;
        RECT 153.400 48.100 153.800 48.200 ;
        RECT 169.400 48.100 169.800 48.200 ;
        RECT 143.800 47.800 151.300 48.100 ;
        RECT 153.400 47.800 169.800 48.100 ;
        RECT 32.600 47.100 33.000 47.200 ;
        RECT 37.400 47.100 37.800 47.200 ;
        RECT 32.600 46.800 37.800 47.100 ;
        RECT 55.800 47.100 56.100 47.800 ;
        RECT 151.000 47.200 151.300 47.800 ;
        RECT 58.200 47.100 58.600 47.200 ;
        RECT 55.800 46.800 58.600 47.100 ;
        RECT 82.200 47.100 82.600 47.200 ;
        RECT 91.800 47.100 92.200 47.200 ;
        RECT 104.600 47.100 105.000 47.200 ;
        RECT 107.000 47.100 107.400 47.200 ;
        RECT 119.800 47.100 120.200 47.200 ;
        RECT 124.600 47.100 125.000 47.200 ;
        RECT 82.200 46.800 125.000 47.100 ;
        RECT 126.200 47.100 126.600 47.200 ;
        RECT 130.200 47.100 130.600 47.200 ;
        RECT 135.000 47.100 135.400 47.200 ;
        RECT 126.200 46.800 135.400 47.100 ;
        RECT 145.400 46.800 145.800 47.200 ;
        RECT 151.000 46.800 151.400 47.200 ;
        RECT 168.600 47.100 169.000 47.200 ;
        RECT 169.400 47.100 169.800 47.200 ;
        RECT 168.600 46.800 169.800 47.100 ;
        RECT 175.000 46.800 175.400 47.200 ;
        RECT 185.400 46.800 185.800 47.200 ;
        RECT 53.400 46.100 53.800 46.300 ;
        RECT 74.200 46.100 74.600 46.200 ;
        RECT 53.400 45.800 74.600 46.100 ;
        RECT 90.200 46.100 90.600 46.200 ;
        RECT 92.600 46.100 93.000 46.200 ;
        RECT 95.000 46.100 95.400 46.200 ;
        RECT 90.200 45.800 95.400 46.100 ;
        RECT 101.400 46.100 101.800 46.200 ;
        RECT 115.000 46.100 115.400 46.200 ;
        RECT 101.400 45.800 115.400 46.100 ;
        RECT 133.400 46.100 133.800 46.200 ;
        RECT 145.400 46.100 145.700 46.800 ;
        RECT 152.600 46.100 153.000 46.200 ;
        RECT 133.400 45.800 153.000 46.100 ;
        RECT 155.000 46.100 155.400 46.200 ;
        RECT 155.800 46.100 156.200 46.200 ;
        RECT 155.000 45.800 156.200 46.100 ;
        RECT 157.400 46.100 157.800 46.200 ;
        RECT 158.200 46.100 158.600 46.200 ;
        RECT 157.400 45.800 158.600 46.100 ;
        RECT 163.800 46.100 164.200 46.300 ;
        RECT 171.000 46.100 171.400 46.200 ;
        RECT 175.000 46.100 175.300 46.800 ;
        RECT 185.400 46.200 185.700 46.800 ;
        RECT 163.800 45.800 175.300 46.100 ;
        RECT 179.800 46.100 180.200 46.200 ;
        RECT 184.600 46.100 185.000 46.200 ;
        RECT 179.800 45.800 185.000 46.100 ;
        RECT 185.400 45.800 185.800 46.200 ;
        RECT 91.000 45.100 91.400 45.200 ;
        RECT 99.000 45.100 99.400 45.200 ;
        RECT 91.000 44.800 99.400 45.100 ;
        RECT 115.800 45.100 116.200 45.200 ;
        RECT 168.600 45.100 169.000 45.200 ;
        RECT 115.800 44.800 169.000 45.100 ;
        RECT 84.600 44.100 85.000 44.200 ;
        RECT 110.200 44.100 110.600 44.200 ;
        RECT 84.600 43.800 110.600 44.100 ;
        RECT 156.600 44.100 157.000 44.200 ;
        RECT 161.400 44.100 161.800 44.200 ;
        RECT 166.200 44.100 166.600 44.200 ;
        RECT 156.600 43.800 166.600 44.100 ;
        RECT 35.800 43.100 36.200 43.200 ;
        RECT 37.400 43.100 37.800 43.200 ;
        RECT 35.800 42.800 37.800 43.100 ;
        RECT 155.000 43.100 155.400 43.200 ;
        RECT 157.400 43.100 157.800 43.200 ;
        RECT 171.000 43.100 171.400 43.200 ;
        RECT 178.200 43.100 178.600 43.200 ;
        RECT 155.000 42.800 178.600 43.100 ;
        RECT 9.400 40.100 9.800 40.200 ;
        RECT 22.200 40.100 22.600 40.200 ;
        RECT 9.400 39.800 22.600 40.100 ;
        RECT 1.400 39.100 1.800 39.200 ;
        RECT 7.800 39.100 8.200 39.200 ;
        RECT 9.400 39.100 9.800 39.200 ;
        RECT 1.400 38.800 9.800 39.100 ;
        RECT 40.600 39.100 41.000 39.200 ;
        RECT 52.600 39.100 53.000 39.200 ;
        RECT 40.600 38.800 53.000 39.100 ;
        RECT 88.600 39.100 89.000 39.200 ;
        RECT 95.800 39.100 96.200 39.200 ;
        RECT 97.400 39.100 97.800 39.200 ;
        RECT 106.200 39.100 106.600 39.200 ;
        RECT 88.600 38.800 106.600 39.100 ;
        RECT 111.800 37.100 112.200 37.200 ;
        RECT 118.200 37.100 118.600 37.200 ;
        RECT 121.400 37.100 121.800 37.200 ;
        RECT 111.800 36.800 121.800 37.100 ;
        RECT 7.000 35.800 7.400 36.200 ;
        RECT 28.600 36.100 29.000 36.200 ;
        RECT 39.000 36.100 39.400 36.200 ;
        RECT 28.600 35.800 39.400 36.100 ;
        RECT 47.800 36.100 48.200 36.200 ;
        RECT 50.200 36.100 50.600 36.200 ;
        RECT 47.800 35.800 50.600 36.100 ;
        RECT 69.400 35.800 69.800 36.200 ;
        RECT 91.800 35.800 92.200 36.200 ;
        RECT 119.000 35.800 119.400 36.200 ;
        RECT 123.800 35.800 124.200 36.200 ;
        RECT 7.000 35.100 7.300 35.800 ;
        RECT 14.200 35.100 14.600 35.200 ;
        RECT 7.000 34.800 14.600 35.100 ;
        RECT 39.800 35.100 40.200 35.200 ;
        RECT 40.600 35.100 41.000 35.200 ;
        RECT 39.800 34.800 41.000 35.100 ;
        RECT 45.400 35.100 45.800 35.200 ;
        RECT 51.800 35.100 52.200 35.200 ;
        RECT 45.400 34.800 52.200 35.100 ;
        RECT 67.800 35.100 68.200 35.200 ;
        RECT 69.400 35.100 69.700 35.800 ;
        RECT 67.800 34.800 69.700 35.100 ;
        RECT 85.400 35.100 85.800 35.200 ;
        RECT 91.800 35.100 92.100 35.800 ;
        RECT 85.400 34.800 92.100 35.100 ;
        RECT 119.000 35.100 119.300 35.800 ;
        RECT 123.800 35.200 124.100 35.800 ;
        RECT 120.600 35.100 121.000 35.200 ;
        RECT 119.000 34.800 121.000 35.100 ;
        RECT 123.800 34.800 124.200 35.200 ;
        RECT 151.800 35.100 152.200 35.200 ;
        RECT 162.200 35.100 162.600 35.200 ;
        RECT 168.600 35.100 169.000 35.200 ;
        RECT 174.200 35.100 174.600 35.200 ;
        RECT 175.000 35.100 175.400 35.200 ;
        RECT 151.800 34.800 162.600 35.100 ;
        RECT 167.800 34.800 175.400 35.100 ;
        RECT 24.600 34.100 25.000 34.200 ;
        RECT 32.600 34.100 33.000 34.200 ;
        RECT 24.600 33.800 33.000 34.100 ;
        RECT 35.800 34.100 36.200 34.200 ;
        RECT 42.200 34.100 42.600 34.200 ;
        RECT 35.800 33.800 42.600 34.100 ;
        RECT 49.400 34.100 49.800 34.200 ;
        RECT 51.000 34.100 51.400 34.200 ;
        RECT 49.400 33.800 51.400 34.100 ;
        RECT 72.600 34.100 73.000 34.200 ;
        RECT 75.000 34.100 75.400 34.200 ;
        RECT 99.000 34.100 99.400 34.200 ;
        RECT 101.400 34.100 101.800 34.400 ;
        RECT 72.600 34.000 101.800 34.100 ;
        RECT 103.800 34.100 104.200 34.200 ;
        RECT 105.400 34.100 105.800 34.200 ;
        RECT 113.400 34.100 113.800 34.200 ;
        RECT 72.600 33.800 101.700 34.000 ;
        RECT 103.800 33.800 113.800 34.100 ;
        RECT 144.600 34.100 145.000 34.200 ;
        RECT 173.400 34.100 173.800 34.200 ;
        RECT 144.600 33.800 173.800 34.100 ;
        RECT 158.200 33.200 158.500 33.800 ;
        RECT 50.200 33.100 50.600 33.200 ;
        RECT 53.400 33.100 53.800 33.200 ;
        RECT 50.200 32.800 53.800 33.100 ;
        RECT 79.000 33.100 79.400 33.200 ;
        RECT 83.800 33.100 84.200 33.200 ;
        RECT 79.000 32.800 84.200 33.100 ;
        RECT 95.000 33.100 95.400 33.200 ;
        RECT 103.800 33.100 104.200 33.200 ;
        RECT 112.600 33.100 113.000 33.200 ;
        RECT 95.000 32.800 113.000 33.100 ;
        RECT 158.200 32.800 158.600 33.200 ;
        RECT 30.200 32.100 30.600 32.200 ;
        RECT 39.800 32.100 40.200 32.200 ;
        RECT 30.200 31.800 40.200 32.100 ;
        RECT 38.200 31.100 38.600 31.200 ;
        RECT 43.000 31.100 43.400 31.200 ;
        RECT 38.200 30.800 43.400 31.100 ;
        RECT 108.600 31.100 109.000 31.200 ;
        RECT 120.600 31.100 121.000 31.200 ;
        RECT 123.800 31.100 124.200 31.200 ;
        RECT 129.400 31.100 129.800 31.200 ;
        RECT 135.000 31.100 135.400 31.200 ;
        RECT 108.600 30.800 135.400 31.100 ;
        RECT 6.200 30.100 6.600 30.200 ;
        RECT 11.000 30.100 11.400 30.200 ;
        RECT 6.200 29.800 11.400 30.100 ;
        RECT 167.800 30.100 168.200 30.200 ;
        RECT 170.200 30.100 170.600 30.200 ;
        RECT 167.800 29.800 170.600 30.100 ;
        RECT 35.000 29.100 35.400 29.200 ;
        RECT 39.800 29.100 40.200 29.200 ;
        RECT 47.800 29.100 48.200 29.200 ;
        RECT 35.000 28.800 36.900 29.100 ;
        RECT 39.800 28.800 48.200 29.100 ;
        RECT 155.000 29.100 155.400 29.200 ;
        RECT 162.200 29.100 162.600 29.200 ;
        RECT 155.000 28.800 162.600 29.100 ;
        RECT 165.400 29.100 165.800 29.200 ;
        RECT 167.000 29.100 167.400 29.200 ;
        RECT 165.400 28.800 167.400 29.100 ;
        RECT 177.400 28.800 177.800 29.200 ;
        RECT 179.000 29.100 179.400 29.200 ;
        RECT 182.200 29.100 182.600 29.200 ;
        RECT 179.000 28.800 182.600 29.100 ;
        RECT 36.600 28.200 36.900 28.800 ;
        RECT 28.600 27.800 29.000 28.200 ;
        RECT 36.600 27.800 37.000 28.200 ;
        RECT 40.600 27.800 41.000 28.200 ;
        RECT 95.800 27.800 96.200 28.200 ;
        RECT 167.000 28.100 167.400 28.200 ;
        RECT 168.600 28.100 169.000 28.200 ;
        RECT 177.400 28.100 177.700 28.800 ;
        RECT 167.000 27.800 177.700 28.100 ;
        RECT 14.200 27.100 14.600 27.200 ;
        RECT 28.600 27.100 28.900 27.800 ;
        RECT 40.600 27.100 40.900 27.800 ;
        RECT 14.200 26.800 40.900 27.100 ;
        RECT 91.800 27.100 92.200 27.200 ;
        RECT 95.800 27.100 96.100 27.800 ;
        RECT 105.400 27.100 105.800 27.200 ;
        RECT 91.800 26.800 105.800 27.100 ;
        RECT 12.600 26.100 13.000 26.200 ;
        RECT 38.200 26.100 38.600 26.200 ;
        RECT 39.800 26.100 40.200 26.200 ;
        RECT 12.600 25.800 20.900 26.100 ;
        RECT 38.200 25.800 40.200 26.100 ;
        RECT 75.000 26.100 75.400 26.200 ;
        RECT 77.400 26.100 77.800 26.200 ;
        RECT 75.000 25.800 77.800 26.100 ;
        RECT 123.800 26.100 124.200 26.200 ;
        RECT 149.400 26.100 149.800 26.200 ;
        RECT 159.800 26.100 160.200 26.200 ;
        RECT 171.800 26.100 172.200 26.200 ;
        RECT 180.600 26.100 181.000 26.200 ;
        RECT 123.800 25.800 133.700 26.100 ;
        RECT 149.400 25.800 157.700 26.100 ;
        RECT 159.800 25.800 181.000 26.100 ;
        RECT 12.600 25.200 12.900 25.800 ;
        RECT 20.600 25.200 20.900 25.800 ;
        RECT 12.600 24.800 13.000 25.200 ;
        RECT 20.600 24.800 21.000 25.200 ;
        RECT 67.800 25.100 68.200 25.200 ;
        RECT 69.400 25.100 69.800 25.200 ;
        RECT 123.800 25.100 124.100 25.800 ;
        RECT 67.800 24.800 124.100 25.100 ;
        RECT 133.400 25.200 133.700 25.800 ;
        RECT 157.400 25.200 157.700 25.800 ;
        RECT 133.400 24.800 133.800 25.200 ;
        RECT 157.400 24.800 157.800 25.200 ;
        RECT 7.800 24.100 8.200 24.200 ;
        RECT 51.000 24.100 51.400 24.200 ;
        RECT 73.400 24.100 73.800 24.200 ;
        RECT 7.800 23.800 73.800 24.100 ;
        RECT 75.800 24.100 76.200 24.200 ;
        RECT 78.200 24.100 78.600 24.200 ;
        RECT 75.800 23.800 78.600 24.100 ;
        RECT 81.400 24.100 81.800 24.200 ;
        RECT 137.400 24.100 137.800 24.200 ;
        RECT 145.400 24.100 145.800 24.200 ;
        RECT 81.400 23.800 145.800 24.100 ;
        RECT 25.400 23.100 25.800 23.200 ;
        RECT 30.200 23.100 30.600 23.200 ;
        RECT 40.600 23.100 41.000 23.200 ;
        RECT 25.400 22.800 41.000 23.100 ;
        RECT 71.800 23.100 72.200 23.200 ;
        RECT 74.200 23.100 74.600 23.200 ;
        RECT 71.800 22.800 74.600 23.100 ;
        RECT 18.200 22.100 18.600 22.200 ;
        RECT 26.200 22.100 26.600 22.200 ;
        RECT 18.200 21.800 26.600 22.100 ;
        RECT 79.000 22.100 79.400 22.200 ;
        RECT 80.600 22.100 81.000 22.200 ;
        RECT 87.000 22.100 87.400 22.200 ;
        RECT 79.000 21.800 87.400 22.100 ;
        RECT 91.800 22.100 92.200 22.200 ;
        RECT 148.600 22.100 149.000 22.200 ;
        RECT 91.800 21.800 149.000 22.100 ;
        RECT 102.200 21.100 102.600 21.200 ;
        RECT 111.800 21.100 112.200 21.200 ;
        RECT 102.200 20.800 112.200 21.100 ;
        RECT 108.600 20.100 109.000 20.200 ;
        RECT 111.000 20.100 111.400 20.200 ;
        RECT 117.400 20.100 117.800 20.200 ;
        RECT 108.600 19.800 117.800 20.100 ;
        RECT 84.600 19.100 85.000 19.200 ;
        RECT 93.400 19.100 93.800 19.200 ;
        RECT 84.600 18.800 93.800 19.100 ;
        RECT 143.000 19.100 143.400 19.200 ;
        RECT 151.800 19.100 152.200 19.200 ;
        RECT 143.000 18.800 152.200 19.100 ;
        RECT 173.400 19.100 173.800 19.200 ;
        RECT 177.400 19.100 177.800 19.200 ;
        RECT 173.400 18.800 177.800 19.100 ;
        RECT 87.800 18.200 88.100 18.800 ;
        RECT 75.800 17.800 76.200 18.200 ;
        RECT 87.800 17.800 88.200 18.200 ;
        RECT 20.600 17.100 21.000 17.200 ;
        RECT 23.800 17.100 24.200 17.200 ;
        RECT 20.600 16.800 24.200 17.100 ;
        RECT 47.000 17.100 47.400 17.200 ;
        RECT 48.600 17.100 49.000 17.200 ;
        RECT 47.000 16.800 49.000 17.100 ;
        RECT 69.400 17.100 69.800 17.200 ;
        RECT 75.800 17.100 76.100 17.800 ;
        RECT 69.400 16.800 76.100 17.100 ;
        RECT 11.000 16.100 11.400 16.200 ;
        RECT 41.400 16.100 41.800 16.200 ;
        RECT 11.000 15.800 41.800 16.100 ;
        RECT 59.800 16.100 60.200 16.200 ;
        RECT 67.000 16.100 67.400 16.200 ;
        RECT 59.800 15.800 67.400 16.100 ;
        RECT 75.000 16.100 75.400 16.200 ;
        RECT 77.400 16.100 77.800 16.200 ;
        RECT 75.000 15.800 77.800 16.100 ;
        RECT 79.000 16.100 79.400 16.200 ;
        RECT 81.400 16.100 81.800 16.200 ;
        RECT 79.000 15.800 81.800 16.100 ;
        RECT 127.800 15.800 128.200 16.200 ;
        RECT 134.200 16.100 134.600 16.200 ;
        RECT 139.800 16.100 140.200 16.200 ;
        RECT 154.200 16.100 154.600 16.200 ;
        RECT 134.200 15.800 154.600 16.100 ;
        RECT 176.600 16.100 177.000 16.200 ;
        RECT 179.800 16.100 180.200 16.200 ;
        RECT 188.600 16.100 189.000 16.200 ;
        RECT 176.600 15.800 189.000 16.100 ;
        RECT 8.600 15.100 9.000 15.200 ;
        RECT 19.000 15.100 19.400 15.200 ;
        RECT 23.800 15.100 24.200 15.200 ;
        RECT 8.600 14.800 17.700 15.100 ;
        RECT 19.000 14.800 24.200 15.100 ;
        RECT 29.400 15.100 29.800 15.200 ;
        RECT 31.800 15.100 32.200 15.200 ;
        RECT 35.000 15.100 35.400 15.200 ;
        RECT 29.400 14.800 35.400 15.100 ;
        RECT 55.800 15.100 56.200 15.200 ;
        RECT 88.600 15.100 89.000 15.200 ;
        RECT 109.400 15.100 109.800 15.200 ;
        RECT 110.200 15.100 110.600 15.200 ;
        RECT 125.400 15.100 125.800 15.200 ;
        RECT 55.800 14.800 125.800 15.100 ;
        RECT 127.800 15.100 128.100 15.800 ;
        RECT 131.800 15.100 132.200 15.200 ;
        RECT 127.800 14.800 132.200 15.100 ;
        RECT 136.600 14.800 137.000 15.200 ;
        RECT 141.400 15.100 141.800 15.200 ;
        RECT 143.800 15.100 144.200 15.200 ;
        RECT 141.400 14.800 144.200 15.100 ;
        RECT 155.000 15.100 155.400 15.200 ;
        RECT 155.800 15.100 156.200 15.200 ;
        RECT 155.000 14.800 156.200 15.100 ;
        RECT 168.600 15.100 169.000 15.200 ;
        RECT 172.600 15.100 173.000 15.200 ;
        RECT 168.600 14.800 173.000 15.100 ;
        RECT 183.800 15.100 184.200 15.200 ;
        RECT 187.800 15.100 188.200 15.200 ;
        RECT 183.800 14.800 188.200 15.100 ;
        RECT 17.400 14.200 17.700 14.800 ;
        RECT 17.400 13.800 17.800 14.200 ;
        RECT 26.200 13.800 26.600 14.200 ;
        RECT 28.600 13.800 29.000 14.200 ;
        RECT 59.800 14.100 60.200 14.200 ;
        RECT 57.400 13.800 60.200 14.100 ;
        RECT 81.400 14.100 81.800 14.200 ;
        RECT 83.800 14.100 84.200 14.200 ;
        RECT 81.400 13.800 84.200 14.100 ;
        RECT 87.000 14.100 87.400 14.200 ;
        RECT 91.800 14.100 92.200 14.200 ;
        RECT 87.000 13.800 92.200 14.100 ;
        RECT 100.600 14.100 101.000 14.200 ;
        RECT 107.800 14.100 108.200 14.200 ;
        RECT 114.200 14.100 114.600 14.200 ;
        RECT 100.600 13.800 114.600 14.100 ;
        RECT 119.000 14.100 119.400 14.200 ;
        RECT 131.000 14.100 131.400 14.200 ;
        RECT 136.600 14.100 136.900 14.800 ;
        RECT 119.000 13.800 136.900 14.100 ;
        RECT 139.000 14.100 139.400 14.200 ;
        RECT 142.200 14.100 142.600 14.200 ;
        RECT 139.000 13.800 142.600 14.100 ;
        RECT 155.000 14.100 155.400 14.200 ;
        RECT 164.600 14.100 165.000 14.200 ;
        RECT 169.400 14.100 169.800 14.200 ;
        RECT 178.200 14.100 178.600 14.200 ;
        RECT 155.000 13.800 178.600 14.100 ;
        RECT 183.000 14.100 183.400 14.200 ;
        RECT 183.800 14.100 184.200 14.200 ;
        RECT 183.000 13.800 184.200 14.100 ;
        RECT 26.200 13.100 26.500 13.800 ;
        RECT 28.600 13.100 28.900 13.800 ;
        RECT 57.400 13.200 57.700 13.800 ;
        RECT 26.200 12.800 28.900 13.100 ;
        RECT 43.000 13.100 43.400 13.200 ;
        RECT 57.400 13.100 57.800 13.200 ;
        RECT 43.000 12.800 57.800 13.100 ;
        RECT 61.400 13.100 61.800 13.200 ;
        RECT 78.200 13.100 78.600 13.200 ;
        RECT 82.200 13.100 82.600 13.200 ;
        RECT 92.600 13.100 93.000 13.200 ;
        RECT 154.200 13.100 154.600 13.200 ;
        RECT 181.400 13.100 181.800 13.200 ;
        RECT 194.200 13.100 194.600 13.200 ;
        RECT 61.400 12.800 181.800 13.100 ;
        RECT 183.000 12.800 194.600 13.100 ;
        RECT 183.000 12.200 183.300 12.800 ;
        RECT 0.600 12.100 1.000 12.200 ;
        RECT 3.800 12.100 4.200 12.200 ;
        RECT 14.200 12.100 14.600 12.200 ;
        RECT 23.000 12.100 23.400 12.200 ;
        RECT 27.000 12.100 27.400 12.200 ;
        RECT 30.200 12.100 30.600 12.200 ;
        RECT 0.600 11.800 30.600 12.100 ;
        RECT 41.400 12.100 41.800 12.200 ;
        RECT 50.200 12.100 50.600 12.200 ;
        RECT 55.000 12.100 55.400 12.200 ;
        RECT 41.400 11.800 55.400 12.100 ;
        RECT 79.000 12.100 79.400 12.200 ;
        RECT 81.400 12.100 81.800 12.200 ;
        RECT 79.000 11.800 81.800 12.100 ;
        RECT 82.200 12.100 82.600 12.200 ;
        RECT 90.200 12.100 90.600 12.200 ;
        RECT 99.000 12.100 99.400 12.200 ;
        RECT 82.200 11.800 99.400 12.100 ;
        RECT 100.600 12.100 101.000 12.200 ;
        RECT 104.600 12.100 105.000 12.200 ;
        RECT 120.600 12.100 121.000 12.200 ;
        RECT 135.800 12.100 136.200 12.200 ;
        RECT 140.600 12.100 141.000 12.200 ;
        RECT 100.600 11.800 105.700 12.100 ;
        RECT 120.600 11.800 141.000 12.100 ;
        RECT 158.200 12.100 158.600 12.200 ;
        RECT 162.200 12.100 162.600 12.200 ;
        RECT 158.200 11.800 162.600 12.100 ;
        RECT 167.000 12.100 167.400 12.200 ;
        RECT 170.200 12.100 170.600 12.200 ;
        RECT 172.600 12.100 173.000 12.200 ;
        RECT 167.000 11.800 173.000 12.100 ;
        RECT 177.400 12.100 177.800 12.200 ;
        RECT 180.600 12.100 181.000 12.200 ;
        RECT 183.000 12.100 183.400 12.200 ;
        RECT 177.400 11.800 183.400 12.100 ;
        RECT 7.000 11.100 7.400 11.200 ;
        RECT 13.400 11.100 13.800 11.200 ;
        RECT 7.000 10.800 13.800 11.100 ;
        RECT 30.200 11.100 30.600 11.200 ;
        RECT 45.400 11.100 45.800 11.200 ;
        RECT 46.200 11.100 46.600 11.200 ;
        RECT 30.200 10.800 46.600 11.100 ;
        RECT 63.800 11.100 64.200 11.200 ;
        RECT 79.000 11.100 79.400 11.200 ;
        RECT 63.800 10.800 79.400 11.100 ;
        RECT 79.800 11.100 80.200 11.200 ;
        RECT 82.200 11.100 82.600 11.200 ;
        RECT 79.800 10.800 82.600 11.100 ;
        RECT 103.800 11.100 104.200 11.200 ;
        RECT 105.400 11.100 105.800 11.200 ;
        RECT 103.800 10.800 105.800 11.100 ;
        RECT 106.200 11.100 106.600 11.200 ;
        RECT 115.000 11.100 115.400 11.200 ;
        RECT 139.800 11.100 140.200 11.200 ;
        RECT 106.200 10.800 140.200 11.100 ;
        RECT 11.800 10.100 12.200 10.200 ;
        RECT 12.600 10.100 13.000 10.200 ;
        RECT 27.000 10.100 27.400 10.200 ;
        RECT 11.800 9.800 27.400 10.100 ;
        RECT 41.400 10.100 41.800 10.200 ;
        RECT 62.200 10.100 62.600 10.200 ;
        RECT 67.000 10.100 67.400 10.200 ;
        RECT 41.400 9.800 67.400 10.100 ;
        RECT 81.400 10.100 81.800 10.200 ;
        RECT 86.200 10.100 86.600 10.200 ;
        RECT 81.400 9.800 86.600 10.100 ;
        RECT 115.800 10.100 116.200 10.200 ;
        RECT 120.600 10.100 121.000 10.200 ;
        RECT 115.800 9.800 121.000 10.100 ;
        RECT 135.000 10.100 135.400 10.200 ;
        RECT 137.400 10.100 137.800 10.200 ;
        RECT 139.000 10.100 139.400 10.200 ;
        RECT 150.200 10.100 150.600 10.200 ;
        RECT 135.000 9.800 136.900 10.100 ;
        RECT 137.400 9.800 150.600 10.100 ;
        RECT 136.600 9.200 136.900 9.800 ;
        RECT 12.600 9.100 13.000 9.200 ;
        RECT 11.800 8.800 13.000 9.100 ;
        RECT 21.400 9.100 21.800 9.200 ;
        RECT 31.000 9.100 31.400 9.200 ;
        RECT 21.400 8.800 31.400 9.100 ;
        RECT 35.800 9.100 36.200 9.200 ;
        RECT 47.000 9.100 47.400 9.200 ;
        RECT 35.800 8.800 47.400 9.100 ;
        RECT 60.600 8.800 61.000 9.200 ;
        RECT 75.000 8.800 75.400 9.200 ;
        RECT 79.000 9.100 79.400 9.200 ;
        RECT 86.200 9.100 86.600 9.200 ;
        RECT 79.000 8.800 86.600 9.100 ;
        RECT 91.800 8.800 92.200 9.200 ;
        RECT 100.600 9.100 101.000 9.200 ;
        RECT 103.800 9.100 104.200 9.200 ;
        RECT 100.600 8.800 104.200 9.100 ;
        RECT 121.400 8.800 121.800 9.200 ;
        RECT 123.000 9.100 123.400 9.200 ;
        RECT 126.200 9.100 126.600 9.200 ;
        RECT 136.600 9.100 137.000 9.200 ;
        RECT 123.000 8.800 137.000 9.100 ;
        RECT 141.400 9.100 141.800 9.200 ;
        RECT 144.600 9.100 145.000 9.200 ;
        RECT 158.200 9.100 158.600 9.200 ;
        RECT 141.400 8.800 158.600 9.100 ;
        RECT 162.200 9.100 162.600 9.200 ;
        RECT 167.000 9.100 167.400 9.200 ;
        RECT 175.800 9.100 176.200 9.200 ;
        RECT 162.200 8.800 176.200 9.100 ;
        RECT 12.600 8.100 13.000 8.200 ;
        RECT 13.400 8.100 13.800 8.200 ;
        RECT 12.600 7.800 13.800 8.100 ;
        RECT 16.600 8.100 17.000 8.200 ;
        RECT 20.600 8.100 21.000 8.200 ;
        RECT 16.600 7.800 21.000 8.100 ;
        RECT 23.800 8.100 24.200 8.200 ;
        RECT 29.400 8.100 29.800 8.200 ;
        RECT 32.600 8.100 33.000 8.200 ;
        RECT 23.800 7.800 33.000 8.100 ;
        RECT 33.400 8.100 33.800 8.200 ;
        RECT 48.600 8.100 49.000 8.200 ;
        RECT 60.600 8.100 60.900 8.800 ;
        RECT 33.400 7.800 60.900 8.100 ;
        RECT 75.000 8.100 75.300 8.800 ;
        RECT 91.800 8.200 92.100 8.800 ;
        RECT 79.800 8.100 80.200 8.200 ;
        RECT 75.000 7.800 80.200 8.100 ;
        RECT 88.600 7.800 89.000 8.200 ;
        RECT 91.800 7.800 92.200 8.200 ;
        RECT 92.600 8.100 93.000 8.200 ;
        RECT 115.000 8.100 115.400 8.200 ;
        RECT 121.400 8.100 121.700 8.800 ;
        RECT 92.600 7.800 121.700 8.100 ;
        RECT 123.000 8.100 123.400 8.200 ;
        RECT 124.600 8.100 125.000 8.200 ;
        RECT 123.000 7.800 125.000 8.100 ;
        RECT 129.400 8.100 129.800 8.200 ;
        RECT 145.400 8.100 145.800 8.200 ;
        RECT 129.400 7.800 145.800 8.100 ;
        RECT 163.000 8.100 163.400 8.200 ;
        RECT 171.800 8.100 172.200 8.200 ;
        RECT 178.200 8.100 178.600 8.200 ;
        RECT 163.000 7.800 178.600 8.100 ;
        RECT 185.400 7.800 185.800 8.200 ;
        RECT 11.000 7.100 11.400 7.200 ;
        RECT 11.800 7.100 12.200 7.200 ;
        RECT 11.000 6.800 12.200 7.100 ;
        RECT 15.800 7.100 16.200 7.200 ;
        RECT 17.400 7.100 17.800 7.200 ;
        RECT 23.000 7.100 23.400 7.200 ;
        RECT 15.800 6.800 23.400 7.100 ;
        RECT 34.200 7.100 34.600 7.200 ;
        RECT 51.800 7.100 52.200 7.200 ;
        RECT 59.000 7.100 59.400 7.200 ;
        RECT 61.400 7.100 61.800 7.200 ;
        RECT 34.200 6.800 61.800 7.100 ;
        RECT 77.400 7.100 77.800 7.200 ;
        RECT 79.000 7.100 79.400 7.200 ;
        RECT 77.400 6.800 79.400 7.100 ;
        RECT 85.400 7.100 85.800 7.200 ;
        RECT 87.800 7.100 88.200 7.200 ;
        RECT 88.600 7.100 88.900 7.800 ;
        RECT 99.800 7.100 100.200 7.200 ;
        RECT 85.400 6.800 88.900 7.100 ;
        RECT 89.400 6.800 100.200 7.100 ;
        RECT 100.600 7.100 101.000 7.200 ;
        RECT 101.400 7.100 101.800 7.200 ;
        RECT 100.600 6.800 101.800 7.100 ;
        RECT 102.200 7.100 102.600 7.200 ;
        RECT 103.000 7.100 103.400 7.200 ;
        RECT 102.200 6.800 103.400 7.100 ;
        RECT 107.000 7.100 107.400 7.200 ;
        RECT 111.800 7.100 112.200 7.200 ;
        RECT 107.000 6.800 112.200 7.100 ;
        RECT 113.400 7.100 113.800 7.200 ;
        RECT 129.400 7.100 129.700 7.800 ;
        RECT 113.400 6.800 129.700 7.100 ;
        RECT 159.000 7.100 159.400 7.200 ;
        RECT 175.800 7.100 176.200 7.200 ;
        RECT 185.400 7.100 185.700 7.800 ;
        RECT 159.000 6.800 185.700 7.100 ;
        RECT 3.800 6.100 4.200 6.200 ;
        RECT 15.000 6.100 15.400 6.200 ;
        RECT 16.600 6.100 17.000 6.200 ;
        RECT 59.800 6.100 60.200 6.200 ;
        RECT 63.800 6.100 64.200 6.200 ;
        RECT 89.400 6.100 89.700 6.800 ;
        RECT 3.800 5.800 16.100 6.100 ;
        RECT 16.600 5.800 89.700 6.100 ;
        RECT 98.200 6.100 98.600 6.200 ;
        RECT 104.600 6.100 105.000 6.200 ;
        RECT 108.600 6.100 109.000 6.200 ;
        RECT 119.800 6.100 120.200 6.200 ;
        RECT 123.800 6.100 124.200 6.200 ;
        RECT 127.000 6.100 127.400 6.200 ;
        RECT 98.200 5.800 123.300 6.100 ;
        RECT 123.800 5.800 127.400 6.100 ;
        RECT 127.800 6.100 128.200 6.200 ;
        RECT 139.000 6.100 139.400 6.200 ;
        RECT 127.800 5.800 139.400 6.100 ;
        RECT 157.400 6.100 157.800 6.200 ;
        RECT 163.000 6.100 163.400 6.200 ;
        RECT 167.800 6.100 168.200 6.200 ;
        RECT 157.400 5.800 168.200 6.100 ;
        RECT 178.200 6.100 178.600 6.200 ;
        RECT 178.200 5.800 182.500 6.100 ;
        RECT 123.000 5.200 123.300 5.800 ;
        RECT 182.200 5.200 182.500 5.800 ;
        RECT 4.600 5.100 5.000 5.200 ;
        RECT 5.400 5.100 5.800 5.200 ;
        RECT 4.600 4.800 5.800 5.100 ;
        RECT 14.200 5.100 14.600 5.200 ;
        RECT 15.800 5.100 16.200 5.200 ;
        RECT 14.200 4.800 16.200 5.100 ;
        RECT 17.400 5.100 17.800 5.200 ;
        RECT 19.800 5.100 20.200 5.200 ;
        RECT 33.400 5.100 33.800 5.200 ;
        RECT 17.400 4.800 33.800 5.100 ;
        RECT 41.400 5.100 41.800 5.200 ;
        RECT 42.200 5.100 42.600 5.200 ;
        RECT 41.400 4.800 42.600 5.100 ;
        RECT 49.400 5.100 49.800 5.200 ;
        RECT 51.000 5.100 51.400 5.200 ;
        RECT 49.400 4.800 51.400 5.100 ;
        RECT 51.800 5.100 52.200 5.200 ;
        RECT 55.000 5.100 55.400 5.200 ;
        RECT 51.800 4.800 55.400 5.100 ;
        RECT 85.400 5.100 85.800 5.200 ;
        RECT 87.800 5.100 88.200 5.200 ;
        RECT 118.200 5.100 118.600 5.200 ;
        RECT 122.200 5.100 122.600 5.200 ;
        RECT 85.400 4.800 122.600 5.100 ;
        RECT 123.000 4.800 123.400 5.200 ;
        RECT 126.200 5.100 126.600 5.200 ;
        RECT 133.400 5.100 133.800 5.200 ;
        RECT 126.200 4.800 133.800 5.100 ;
        RECT 182.200 4.800 182.600 5.200 ;
        RECT 25.400 4.100 25.800 4.200 ;
        RECT 29.400 4.100 29.800 4.200 ;
        RECT 53.400 4.100 53.800 4.200 ;
        RECT 84.600 4.100 85.000 4.200 ;
        RECT 25.400 3.800 85.000 4.100 ;
        RECT 103.000 4.100 103.400 4.200 ;
        RECT 107.000 4.100 107.400 4.200 ;
        RECT 103.000 3.800 107.400 4.100 ;
        RECT 122.200 4.100 122.500 4.800 ;
        RECT 163.000 4.100 163.400 4.200 ;
        RECT 122.200 3.800 163.400 4.100 ;
      LAYER via3 ;
        RECT 165.400 161.800 165.800 162.200 ;
        RECT 60.600 153.800 61.000 154.200 ;
        RECT 95.800 152.800 96.200 153.200 ;
        RECT 81.400 150.800 81.800 151.200 ;
        RECT 102.200 147.800 102.600 148.200 ;
        RECT 123.000 145.800 123.400 146.200 ;
        RECT 95.800 144.800 96.200 145.200 ;
        RECT 124.600 144.800 125.000 145.200 ;
        RECT 12.600 143.800 13.000 144.200 ;
        RECT 190.200 142.800 190.600 143.200 ;
        RECT 44.600 138.800 45.000 139.200 ;
        RECT 79.000 137.800 79.400 138.200 ;
        RECT 173.400 137.800 173.800 138.200 ;
        RECT 27.800 135.800 28.200 136.200 ;
        RECT 75.800 134.800 76.200 135.200 ;
        RECT 123.000 134.800 123.400 135.200 ;
        RECT 130.200 134.800 130.600 135.200 ;
        RECT 165.400 134.800 165.800 135.200 ;
        RECT 56.600 133.800 57.000 134.200 ;
        RECT 141.400 133.800 141.800 134.200 ;
        RECT 158.200 133.800 158.600 134.200 ;
        RECT 89.400 130.800 89.800 131.200 ;
        RECT 84.600 129.800 85.000 130.200 ;
        RECT 159.800 126.800 160.200 127.200 ;
        RECT 193.400 126.800 193.800 127.200 ;
        RECT 59.800 125.800 60.200 126.200 ;
        RECT 38.200 124.800 38.600 125.200 ;
        RECT 40.600 124.800 41.000 125.200 ;
        RECT 139.800 124.800 140.200 125.200 ;
        RECT 128.600 122.800 129.000 123.200 ;
        RECT 174.200 121.800 174.600 122.200 ;
        RECT 82.200 119.800 82.600 120.200 ;
        RECT 35.800 114.800 36.200 115.200 ;
        RECT 12.600 113.800 13.000 114.200 ;
        RECT 27.000 113.800 27.400 114.200 ;
        RECT 87.000 113.800 87.400 114.200 ;
        RECT 194.200 112.800 194.600 113.200 ;
        RECT 27.000 108.800 27.400 109.200 ;
        RECT 37.400 108.800 37.800 109.200 ;
        RECT 39.800 107.800 40.200 108.200 ;
        RECT 92.600 107.800 93.000 108.200 ;
        RECT 37.400 106.800 37.800 107.200 ;
        RECT 48.600 105.800 49.000 106.200 ;
        RECT 55.800 101.800 56.200 102.200 ;
        RECT 128.600 98.800 129.000 99.200 ;
        RECT 112.600 97.800 113.000 98.200 ;
        RECT 42.200 96.800 42.600 97.200 ;
        RECT 130.200 95.800 130.600 96.200 ;
        RECT 17.400 94.800 17.800 95.200 ;
        RECT 39.800 94.800 40.200 95.200 ;
        RECT 126.200 94.800 126.600 95.200 ;
        RECT 8.600 93.800 9.000 94.200 ;
        RECT 45.400 93.800 45.800 94.200 ;
        RECT 132.600 91.800 133.000 92.200 ;
        RECT 10.200 90.800 10.600 91.200 ;
        RECT 15.800 90.800 16.200 91.200 ;
        RECT 39.800 89.800 40.200 90.200 ;
        RECT 51.000 89.800 51.400 90.200 ;
        RECT 57.400 88.800 57.800 89.200 ;
        RECT 184.600 88.800 185.000 89.200 ;
        RECT 58.200 87.800 58.600 88.200 ;
        RECT 8.600 85.800 9.000 86.200 ;
        RECT 11.800 85.800 12.200 86.200 ;
        RECT 138.200 85.800 138.600 86.200 ;
        RECT 47.800 84.800 48.200 85.200 ;
        RECT 139.800 83.800 140.200 84.200 ;
        RECT 50.200 81.800 50.600 82.200 ;
        RECT 80.600 81.800 81.000 82.200 ;
        RECT 171.000 81.800 171.400 82.200 ;
        RECT 88.600 79.800 89.000 80.200 ;
        RECT 89.400 77.800 89.800 78.200 ;
        RECT 40.600 75.800 41.000 76.200 ;
        RECT 166.200 74.800 166.600 75.200 ;
        RECT 39.800 73.800 40.200 74.200 ;
        RECT 63.800 72.800 64.200 73.200 ;
        RECT 63.000 68.800 63.400 69.200 ;
        RECT 123.800 67.800 124.200 68.200 ;
        RECT 79.800 66.800 80.200 67.200 ;
        RECT 171.000 65.800 171.400 66.200 ;
        RECT 84.600 63.800 85.000 64.200 ;
        RECT 80.600 57.800 81.000 58.200 ;
        RECT 169.400 57.800 169.800 58.200 ;
        RECT 185.400 56.800 185.800 57.200 ;
        RECT 47.800 54.800 48.200 55.200 ;
        RECT 114.200 54.800 114.600 55.200 ;
        RECT 84.600 53.800 85.000 54.200 ;
        RECT 178.200 53.800 178.600 54.200 ;
        RECT 194.200 52.800 194.600 53.200 ;
        RECT 183.800 48.800 184.200 49.200 ;
        RECT 169.400 46.800 169.800 47.200 ;
        RECT 37.400 42.800 37.800 43.200 ;
        RECT 171.000 42.800 171.400 43.200 ;
        RECT 7.800 38.800 8.200 39.200 ;
        RECT 83.800 32.800 84.200 33.200 ;
        RECT 39.800 31.800 40.200 32.200 ;
        RECT 39.800 25.800 40.200 26.200 ;
        RECT 151.800 18.800 152.200 19.200 ;
        RECT 155.800 14.800 156.200 15.200 ;
        RECT 114.200 13.800 114.600 14.200 ;
        RECT 79.000 10.800 79.400 11.200 ;
        RECT 12.600 8.800 13.000 9.200 ;
        RECT 11.800 6.800 12.200 7.200 ;
        RECT 101.400 6.800 101.800 7.200 ;
        RECT 103.000 6.800 103.400 7.200 ;
        RECT 33.400 4.800 33.800 5.200 ;
        RECT 42.200 4.800 42.600 5.200 ;
      LAYER metal4 ;
        RECT 102.200 163.800 102.600 164.200 ;
        RECT 86.200 161.800 86.600 162.200 ;
        RECT 43.800 158.100 44.200 158.200 ;
        RECT 43.800 157.800 44.900 158.100 ;
        RECT 40.600 146.800 41.000 147.200 ;
        RECT 12.600 143.800 13.000 144.200 ;
        RECT 11.800 134.800 12.200 135.200 ;
        RECT 9.400 117.100 9.800 117.200 ;
        RECT 9.400 116.800 10.500 117.100 ;
        RECT 10.200 96.200 10.500 116.800 ;
        RECT 10.200 95.800 10.600 96.200 ;
        RECT 8.600 94.100 9.000 94.200 ;
        RECT 7.800 93.800 9.000 94.100 ;
        RECT 7.800 92.200 8.100 93.800 ;
        RECT 7.800 91.800 8.200 92.200 ;
        RECT 7.800 39.200 8.100 91.800 ;
        RECT 10.200 91.200 10.500 95.800 ;
        RECT 10.200 90.800 10.600 91.200 ;
        RECT 11.800 86.200 12.100 134.800 ;
        RECT 12.600 114.200 12.900 143.800 ;
        RECT 27.800 136.100 28.200 136.200 ;
        RECT 27.000 135.800 28.200 136.100 ;
        RECT 37.400 135.800 37.800 136.200 ;
        RECT 27.000 127.200 27.300 135.800 ;
        RECT 27.000 126.800 27.400 127.200 ;
        RECT 15.000 126.100 15.400 126.200 ;
        RECT 15.000 125.800 16.100 126.100 ;
        RECT 12.600 113.800 13.000 114.200 ;
        RECT 12.600 107.200 12.900 113.800 ;
        RECT 12.600 106.800 13.000 107.200 ;
        RECT 15.800 91.200 16.100 125.800 ;
        RECT 27.000 114.200 27.300 126.800 ;
        RECT 37.400 125.100 37.700 135.800 ;
        RECT 40.600 125.200 40.900 146.800 ;
        RECT 44.600 139.200 44.900 157.800 ;
        RECT 60.600 153.800 61.000 154.200 ;
        RECT 44.600 138.800 45.000 139.200 ;
        RECT 56.600 134.100 57.000 134.200 ;
        RECT 55.800 133.800 57.000 134.100 ;
        RECT 38.200 125.100 38.600 125.200 ;
        RECT 37.400 124.800 38.600 125.100 ;
        RECT 40.600 124.800 41.000 125.200 ;
        RECT 35.800 114.800 36.200 115.200 ;
        RECT 27.000 113.800 27.400 114.200 ;
        RECT 27.000 109.200 27.300 113.800 ;
        RECT 27.000 108.800 27.400 109.200 ;
        RECT 35.800 103.200 36.100 114.800 ;
        RECT 37.400 108.800 37.800 109.200 ;
        RECT 37.400 107.200 37.700 108.800 ;
        RECT 39.800 108.100 40.200 108.200 ;
        RECT 40.600 108.100 40.900 124.800 ;
        RECT 39.800 107.800 40.900 108.100 ;
        RECT 47.800 120.800 48.200 121.200 ;
        RECT 37.400 106.800 37.800 107.200 ;
        RECT 47.800 106.100 48.100 120.800 ;
        RECT 50.200 106.800 50.600 107.200 ;
        RECT 48.600 106.100 49.000 106.200 ;
        RECT 47.800 105.800 49.000 106.100 ;
        RECT 35.800 102.800 36.200 103.200 ;
        RECT 42.200 96.800 42.600 97.200 ;
        RECT 43.800 96.800 44.200 97.200 ;
        RECT 40.600 95.800 41.000 96.200 ;
        RECT 17.400 95.100 17.800 95.200 ;
        RECT 18.200 95.100 18.600 95.200 ;
        RECT 17.400 94.800 18.600 95.100 ;
        RECT 39.000 95.100 39.400 95.200 ;
        RECT 39.800 95.100 40.200 95.200 ;
        RECT 39.000 94.800 40.200 95.100 ;
        RECT 25.400 94.100 25.800 94.200 ;
        RECT 26.200 94.100 26.600 94.200 ;
        RECT 25.400 93.800 26.600 94.100 ;
        RECT 15.800 90.800 16.200 91.200 ;
        RECT 39.800 89.800 40.200 90.200 ;
        RECT 37.400 88.800 37.800 89.200 ;
        RECT 8.600 85.800 9.000 86.200 ;
        RECT 11.800 85.800 12.200 86.200 ;
        RECT 8.600 56.200 8.900 85.800 ;
        RECT 8.600 55.800 9.000 56.200 ;
        RECT 37.400 43.200 37.700 88.800 ;
        RECT 39.800 79.200 40.100 89.800 ;
        RECT 38.200 78.800 38.600 79.200 ;
        RECT 39.800 78.800 40.200 79.200 ;
        RECT 38.200 49.200 38.500 78.800 ;
        RECT 40.600 76.200 40.900 95.800 ;
        RECT 42.200 95.200 42.500 96.800 ;
        RECT 41.400 94.800 41.800 95.200 ;
        RECT 42.200 94.800 42.600 95.200 ;
        RECT 41.400 94.200 41.700 94.800 ;
        RECT 41.400 93.800 41.800 94.200 ;
        RECT 43.800 87.200 44.100 96.800 ;
        RECT 45.400 93.800 45.800 94.200 ;
        RECT 45.400 91.200 45.700 93.800 ;
        RECT 45.400 90.800 45.800 91.200 ;
        RECT 43.800 86.800 44.200 87.200 ;
        RECT 47.800 84.800 48.200 85.200 ;
        RECT 40.600 75.800 41.000 76.200 ;
        RECT 39.800 73.800 40.200 74.200 ;
        RECT 38.200 48.800 38.600 49.200 ;
        RECT 37.400 42.800 37.800 43.200 ;
        RECT 7.800 38.800 8.200 39.200 ;
        RECT 39.800 35.200 40.100 73.800 ;
        RECT 47.800 65.200 48.100 84.800 ;
        RECT 50.200 82.200 50.500 106.800 ;
        RECT 55.800 102.200 56.100 133.800 ;
        RECT 59.800 125.800 60.200 126.200 ;
        RECT 59.800 124.200 60.100 125.800 ;
        RECT 59.800 123.800 60.200 124.200 ;
        RECT 57.400 122.800 57.800 123.200 ;
        RECT 55.800 101.800 56.200 102.200 ;
        RECT 51.000 91.800 51.400 92.200 ;
        RECT 51.000 90.200 51.300 91.800 ;
        RECT 51.000 89.800 51.400 90.200 ;
        RECT 57.400 89.200 57.700 122.800 ;
        RECT 59.800 114.800 60.200 115.200 ;
        RECT 58.200 93.800 58.600 94.200 ;
        RECT 57.400 88.800 57.800 89.200 ;
        RECT 58.200 88.200 58.500 93.800 ;
        RECT 58.200 87.800 58.600 88.200 ;
        RECT 59.800 86.200 60.100 114.800 ;
        RECT 60.600 110.200 60.900 153.800 ;
        RECT 81.400 151.100 81.800 151.200 ;
        RECT 80.600 150.800 81.800 151.100 ;
        RECT 79.000 137.800 79.400 138.200 ;
        RECT 73.400 136.800 73.800 137.200 ;
        RECT 73.400 125.200 73.700 136.800 ;
        RECT 75.800 134.800 76.200 135.200 ;
        RECT 75.800 133.200 76.100 134.800 ;
        RECT 75.800 132.800 76.200 133.200 ;
        RECT 73.400 124.800 73.800 125.200 ;
        RECT 60.600 109.800 61.000 110.200 ;
        RECT 59.800 85.800 60.200 86.200 ;
        RECT 50.200 81.800 50.600 82.200 ;
        RECT 78.200 75.800 78.600 76.200 ;
        RECT 77.400 74.800 77.800 75.200 ;
        RECT 63.800 73.800 64.200 74.200 ;
        RECT 63.800 73.200 64.100 73.800 ;
        RECT 63.800 72.800 64.200 73.200 ;
        RECT 63.000 70.800 63.400 71.200 ;
        RECT 63.000 69.200 63.300 70.800 ;
        RECT 77.400 69.200 77.700 74.800 ;
        RECT 78.200 73.200 78.500 75.800 ;
        RECT 78.200 72.800 78.600 73.200 ;
        RECT 63.000 68.800 63.400 69.200 ;
        RECT 77.400 68.800 77.800 69.200 ;
        RECT 47.800 64.800 48.200 65.200 ;
        RECT 47.800 56.800 48.200 57.200 ;
        RECT 47.800 55.200 48.100 56.800 ;
        RECT 47.800 54.800 48.200 55.200 ;
        RECT 79.000 50.200 79.300 137.800 ;
        RECT 80.600 128.200 80.900 150.800 ;
        RECT 84.600 129.800 85.000 130.200 ;
        RECT 80.600 127.800 81.000 128.200 ;
        RECT 82.200 120.100 82.600 120.200 ;
        RECT 81.400 119.800 82.600 120.100 ;
        RECT 79.800 110.800 80.200 111.200 ;
        RECT 79.800 75.200 80.100 110.800 ;
        RECT 81.400 106.200 81.700 119.800 ;
        RECT 81.400 105.800 81.800 106.200 ;
        RECT 80.600 81.800 81.000 82.200 ;
        RECT 79.800 74.800 80.200 75.200 ;
        RECT 79.800 67.200 80.100 74.800 ;
        RECT 79.800 66.800 80.200 67.200 ;
        RECT 80.600 58.200 80.900 81.800 ;
        RECT 84.600 75.200 84.900 129.800 ;
        RECT 86.200 114.100 86.500 161.800 ;
        RECT 95.800 152.800 96.200 153.200 ;
        RECT 95.800 145.200 96.100 152.800 ;
        RECT 102.200 148.200 102.500 163.800 ;
        RECT 124.600 161.800 125.000 162.200 ;
        RECT 165.400 161.800 165.800 162.200 ;
        RECT 102.200 147.800 102.600 148.200 ;
        RECT 123.000 147.800 123.400 148.200 ;
        RECT 123.000 146.200 123.300 147.800 ;
        RECT 123.000 145.800 123.400 146.200 ;
        RECT 124.600 145.200 124.900 161.800 ;
        RECT 165.400 153.200 165.700 161.800 ;
        RECT 174.200 154.800 174.600 155.200 ;
        RECT 165.400 152.800 165.800 153.200 ;
        RECT 162.200 147.800 162.600 148.200 ;
        RECT 162.200 145.200 162.500 147.800 ;
        RECT 95.800 144.800 96.200 145.200 ;
        RECT 124.600 144.800 125.000 145.200 ;
        RECT 162.200 144.800 162.600 145.200 ;
        RECT 138.200 142.800 138.600 143.200 ;
        RECT 111.800 137.800 112.200 138.200 ;
        RECT 92.600 134.800 93.000 135.200 ;
        RECT 89.400 130.800 89.800 131.200 ;
        RECT 87.000 114.100 87.400 114.200 ;
        RECT 86.200 113.800 87.400 114.100 ;
        RECT 88.600 79.800 89.000 80.200 ;
        RECT 84.600 74.800 85.000 75.200 ;
        RECT 84.600 64.200 84.900 74.800 ;
        RECT 84.600 63.800 85.000 64.200 ;
        RECT 80.600 57.800 81.000 58.200 ;
        RECT 80.600 57.200 80.900 57.800 ;
        RECT 80.600 56.800 81.000 57.200 ;
        RECT 84.600 54.100 85.000 54.200 ;
        RECT 83.800 53.800 85.000 54.100 ;
        RECT 83.800 52.200 84.100 53.800 ;
        RECT 83.800 51.800 84.200 52.200 ;
        RECT 79.000 49.800 79.400 50.200 ;
        RECT 67.800 47.800 68.200 48.200 ;
        RECT 39.800 34.800 40.200 35.200 ;
        RECT 39.800 32.200 40.100 34.800 ;
        RECT 39.800 31.800 40.200 32.200 ;
        RECT 39.800 29.200 40.100 31.800 ;
        RECT 39.800 28.800 40.200 29.200 ;
        RECT 39.800 26.200 40.100 28.800 ;
        RECT 39.800 25.800 40.200 26.200 ;
        RECT 67.800 25.200 68.100 47.800 ;
        RECT 83.800 33.200 84.100 51.800 ;
        RECT 88.600 49.200 88.900 79.800 ;
        RECT 89.400 78.200 89.700 130.800 ;
        RECT 92.600 108.200 92.900 134.800 ;
        RECT 92.600 107.800 93.000 108.200 ;
        RECT 111.800 98.100 112.100 137.800 ;
        RECT 123.000 134.800 123.400 135.200 ;
        RECT 130.200 134.800 130.600 135.200 ;
        RECT 123.000 112.200 123.300 134.800 ;
        RECT 128.600 122.800 129.000 123.200 ;
        RECT 123.000 111.800 123.400 112.200 ;
        RECT 128.600 99.200 128.900 122.800 ;
        RECT 130.200 115.200 130.500 134.800 ;
        RECT 138.200 124.200 138.500 142.800 ;
        RECT 159.000 138.800 159.400 139.200 ;
        RECT 141.400 134.100 141.800 134.200 ;
        RECT 142.200 134.100 142.600 134.200 ;
        RECT 141.400 133.800 142.600 134.100 ;
        RECT 157.400 134.100 157.800 134.200 ;
        RECT 158.200 134.100 158.600 134.200 ;
        RECT 157.400 133.800 158.600 134.100 ;
        RECT 139.800 124.800 140.200 125.200 ;
        RECT 138.200 123.800 138.600 124.200 ;
        RECT 130.200 114.800 130.600 115.200 ;
        RECT 128.600 98.800 129.000 99.200 ;
        RECT 112.600 98.100 113.000 98.200 ;
        RECT 111.800 97.800 113.000 98.100 ;
        RECT 126.200 95.100 126.600 95.200 ;
        RECT 125.400 94.800 126.600 95.100 ;
        RECT 104.600 88.800 105.000 89.200 ;
        RECT 104.600 86.200 104.900 88.800 ;
        RECT 104.600 85.800 105.000 86.200 ;
        RECT 89.400 77.800 89.800 78.200 ;
        RECT 125.400 75.200 125.700 94.800 ;
        RECT 128.600 94.200 128.900 98.800 ;
        RECT 130.200 96.200 130.500 114.800 ;
        RECT 130.200 95.800 130.600 96.200 ;
        RECT 128.600 93.800 129.000 94.200 ;
        RECT 130.200 91.200 130.500 95.800 ;
        RECT 131.800 92.100 132.200 92.200 ;
        RECT 132.600 92.100 133.000 92.200 ;
        RECT 131.800 91.800 133.000 92.100 ;
        RECT 130.200 90.800 130.600 91.200 ;
        RECT 138.200 86.200 138.500 123.800 ;
        RECT 139.800 119.200 140.100 124.800 ;
        RECT 139.800 118.800 140.200 119.200 ;
        RECT 138.200 85.800 138.600 86.200 ;
        RECT 139.800 84.200 140.100 118.800 ;
        RECT 139.800 83.800 140.200 84.200 ;
        RECT 125.400 74.800 125.800 75.200 ;
        RECT 107.000 72.800 107.400 73.200 ;
        RECT 151.800 72.800 152.200 73.200 ;
        RECT 107.000 66.200 107.300 72.800 ;
        RECT 123.800 67.800 124.200 68.200 ;
        RECT 107.000 65.800 107.400 66.200 ;
        RECT 114.200 54.800 114.600 55.200 ;
        RECT 114.200 54.200 114.500 54.800 ;
        RECT 114.200 53.800 114.600 54.200 ;
        RECT 119.000 54.100 119.400 54.200 ;
        RECT 119.800 54.100 120.200 54.200 ;
        RECT 119.000 53.800 120.200 54.100 ;
        RECT 88.600 48.800 89.000 49.200 ;
        RECT 123.800 35.200 124.100 67.800 ;
        RECT 123.800 34.800 124.200 35.200 ;
        RECT 83.800 32.800 84.200 33.200 ;
        RECT 91.800 26.800 92.200 27.200 ;
        RECT 12.600 24.800 13.000 25.200 ;
        RECT 67.800 24.800 68.200 25.200 ;
        RECT 11.800 9.800 12.200 10.200 ;
        RECT 11.800 7.200 12.100 9.800 ;
        RECT 12.600 9.200 12.900 24.800 ;
        RECT 79.000 15.800 79.400 16.200 ;
        RECT 41.400 11.800 41.800 12.200 ;
        RECT 12.600 8.800 13.000 9.200 ;
        RECT 12.600 8.100 13.000 8.200 ;
        RECT 13.400 8.100 13.800 8.200 ;
        RECT 12.600 7.800 13.800 8.100 ;
        RECT 33.400 7.800 33.800 8.200 ;
        RECT 11.800 6.800 12.200 7.200 ;
        RECT 33.400 5.200 33.700 7.800 ;
        RECT 4.600 5.100 5.000 5.200 ;
        RECT 5.400 5.100 5.800 5.200 ;
        RECT 4.600 4.800 5.800 5.100 ;
        RECT 16.600 5.100 17.000 5.200 ;
        RECT 17.400 5.100 17.800 5.200 ;
        RECT 16.600 4.800 17.800 5.100 ;
        RECT 33.400 4.800 33.800 5.200 ;
        RECT 41.400 5.100 41.700 11.800 ;
        RECT 79.000 11.200 79.300 15.800 ;
        RECT 79.000 10.800 79.400 11.200 ;
        RECT 91.800 8.200 92.100 26.800 ;
        RECT 123.800 26.200 124.100 34.800 ;
        RECT 123.800 25.800 124.200 26.200 ;
        RECT 151.800 19.200 152.100 72.800 ;
        RECT 159.000 66.200 159.300 138.800 ;
        RECT 165.400 135.200 165.700 152.800 ;
        RECT 173.400 137.800 173.800 138.200 ;
        RECT 165.400 134.800 165.800 135.200 ;
        RECT 159.800 126.800 160.200 127.200 ;
        RECT 159.800 89.200 160.100 126.800 ;
        RECT 165.400 124.200 165.700 134.800 ;
        RECT 165.400 123.800 165.800 124.200 ;
        RECT 173.400 106.200 173.700 137.800 ;
        RECT 174.200 122.200 174.500 154.800 ;
        RECT 190.200 142.800 190.600 143.200 ;
        RECT 174.200 121.800 174.600 122.200 ;
        RECT 190.200 106.200 190.500 142.800 ;
        RECT 193.400 126.800 193.800 127.200 ;
        RECT 173.400 105.800 173.800 106.200 ;
        RECT 190.200 105.800 190.600 106.200 ;
        RECT 166.200 94.800 166.600 95.200 ;
        RECT 159.800 88.800 160.200 89.200 ;
        RECT 166.200 75.200 166.500 94.800 ;
        RECT 184.600 88.800 185.000 89.200 ;
        RECT 171.000 81.800 171.400 82.200 ;
        RECT 166.200 74.800 166.600 75.200 ;
        RECT 171.000 73.200 171.300 81.800 ;
        RECT 184.600 74.200 184.900 88.800 ;
        RECT 184.600 73.800 185.000 74.200 ;
        RECT 171.000 72.800 171.400 73.200 ;
        RECT 171.000 66.200 171.300 72.800 ;
        RECT 159.000 65.800 159.400 66.200 ;
        RECT 171.000 65.800 171.400 66.200 ;
        RECT 169.400 57.800 169.800 58.200 ;
        RECT 169.400 47.200 169.700 57.800 ;
        RECT 169.400 46.800 169.800 47.200 ;
        RECT 171.000 43.200 171.300 65.800 ;
        RECT 193.400 59.200 193.700 126.800 ;
        RECT 194.200 112.800 194.600 113.200 ;
        RECT 193.400 58.800 193.800 59.200 ;
        RECT 185.400 56.800 185.800 57.200 ;
        RECT 178.200 53.800 178.600 54.200 ;
        RECT 171.000 42.800 171.400 43.200 ;
        RECT 151.800 18.800 152.200 19.200 ;
        RECT 114.200 14.800 114.600 15.200 ;
        RECT 155.000 15.100 155.400 15.200 ;
        RECT 155.800 15.100 156.200 15.200 ;
        RECT 155.000 14.800 156.200 15.100 ;
        RECT 114.200 14.200 114.500 14.800 ;
        RECT 114.200 13.800 114.600 14.200 ;
        RECT 51.800 7.800 52.200 8.200 ;
        RECT 88.600 7.800 89.000 8.200 ;
        RECT 91.800 7.800 92.200 8.200 ;
        RECT 51.800 5.200 52.100 7.800 ;
        RECT 88.600 7.200 88.900 7.800 ;
        RECT 88.600 6.800 89.000 7.200 ;
        RECT 100.600 7.100 101.000 7.200 ;
        RECT 101.400 7.100 101.800 7.200 ;
        RECT 100.600 6.800 101.800 7.100 ;
        RECT 102.200 7.100 102.600 7.200 ;
        RECT 103.000 7.100 103.400 7.200 ;
        RECT 102.200 6.800 103.400 7.100 ;
        RECT 123.800 6.800 124.200 7.200 ;
        RECT 123.800 6.200 124.100 6.800 ;
        RECT 178.200 6.200 178.500 53.800 ;
        RECT 183.800 48.800 184.200 49.200 ;
        RECT 183.000 14.100 183.400 14.200 ;
        RECT 183.800 14.100 184.100 48.800 ;
        RECT 185.400 46.200 185.700 56.800 ;
        RECT 194.200 53.200 194.500 112.800 ;
        RECT 194.200 52.800 194.600 53.200 ;
        RECT 185.400 45.800 185.800 46.200 ;
        RECT 183.000 13.800 184.100 14.100 ;
        RECT 123.800 5.800 124.200 6.200 ;
        RECT 178.200 5.800 178.600 6.200 ;
        RECT 42.200 5.100 42.600 5.200 ;
        RECT 41.400 4.800 42.600 5.100 ;
        RECT 51.800 4.800 52.200 5.200 ;
      LAYER via4 ;
        RECT 18.200 94.800 18.600 95.200 ;
        RECT 26.200 93.800 26.600 94.200 ;
        RECT 142.200 133.800 142.600 134.200 ;
        RECT 119.800 53.800 120.200 54.200 ;
        RECT 13.400 7.800 13.800 8.200 ;
        RECT 5.400 4.800 5.800 5.200 ;
      LAYER metal5 ;
        RECT 142.200 134.100 142.600 134.200 ;
        RECT 157.400 134.100 157.800 134.200 ;
        RECT 142.200 133.800 157.800 134.100 ;
        RECT 18.200 95.100 18.600 95.200 ;
        RECT 39.000 95.100 39.400 95.200 ;
        RECT 18.200 94.800 39.400 95.100 ;
        RECT 26.200 94.100 26.600 94.200 ;
        RECT 41.400 94.100 41.800 94.200 ;
        RECT 26.200 93.800 41.800 94.100 ;
        RECT 51.000 92.100 51.400 92.200 ;
        RECT 131.800 92.100 132.200 92.200 ;
        RECT 51.000 91.800 132.200 92.100 ;
        RECT 63.800 73.800 64.200 74.200 ;
        RECT 63.800 73.100 64.100 73.800 ;
        RECT 78.200 73.100 78.600 73.200 ;
        RECT 63.800 72.800 78.600 73.100 ;
        RECT 114.200 54.100 114.600 54.200 ;
        RECT 119.800 54.100 120.200 54.200 ;
        RECT 114.200 53.800 120.200 54.100 ;
        RECT 114.200 15.100 114.600 15.200 ;
        RECT 155.000 15.100 155.400 15.200 ;
        RECT 114.200 14.800 155.400 15.100 ;
        RECT 13.400 8.100 13.800 8.200 ;
        RECT 51.800 8.100 52.200 8.200 ;
        RECT 13.400 7.800 52.200 8.100 ;
        RECT 88.600 7.100 89.000 7.200 ;
        RECT 100.600 7.100 101.000 7.200 ;
        RECT 88.600 6.800 101.000 7.100 ;
        RECT 102.200 7.100 102.600 7.200 ;
        RECT 123.800 7.100 124.200 7.200 ;
        RECT 102.200 6.800 124.200 7.100 ;
        RECT 5.400 5.100 5.800 5.200 ;
        RECT 16.600 5.100 17.000 5.200 ;
        RECT 5.400 4.800 17.000 5.100 ;
  END
END alarm_clock_top
END LIBRARY

