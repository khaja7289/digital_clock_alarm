magic
tech scmos
timestamp 1696677024
<< metal1 >>
rect 968 1703 970 1707
rect 974 1703 977 1707
rect 981 1703 984 1707
rect 86 1671 89 1681
rect 1514 1678 1515 1682
rect 86 1668 94 1671
rect 1454 1668 1465 1671
rect 54 1661 57 1668
rect 46 1658 57 1661
rect 190 1658 209 1661
rect 450 1658 465 1661
rect 542 1658 550 1661
rect 614 1658 622 1661
rect 674 1658 689 1661
rect 838 1658 857 1661
rect 890 1658 897 1661
rect 1454 1662 1457 1668
rect 1018 1658 1033 1661
rect 1330 1658 1337 1661
rect 1790 1658 1798 1661
rect 1934 1618 1942 1621
rect 456 1603 458 1607
rect 462 1603 465 1607
rect 469 1603 472 1607
rect 1480 1603 1482 1607
rect 1486 1603 1489 1607
rect 1493 1603 1496 1607
rect 125 1588 126 1592
rect 1122 1588 1123 1592
rect 1674 1588 1675 1592
rect 1813 1588 1814 1592
rect 314 1568 317 1572
rect 826 1568 829 1572
rect 974 1568 982 1571
rect 1603 1568 1606 1572
rect 106 1548 113 1551
rect 1038 1548 1057 1551
rect 1166 1548 1185 1551
rect 1190 1548 1201 1551
rect 1230 1551 1233 1561
rect 1226 1548 1233 1551
rect 1246 1548 1254 1551
rect 1334 1548 1345 1551
rect 1490 1548 1502 1551
rect 1654 1548 1662 1551
rect 1342 1542 1345 1548
rect 154 1538 161 1541
rect 974 1538 1001 1541
rect 1258 1538 1265 1541
rect 1446 1541 1449 1548
rect 1654 1546 1658 1548
rect 1438 1538 1449 1541
rect 1678 1541 1681 1551
rect 1726 1548 1734 1551
rect 1774 1541 1777 1548
rect 1678 1538 1697 1541
rect 1766 1538 1777 1541
rect 1822 1538 1834 1541
rect 1942 1538 1950 1541
rect 974 1532 977 1538
rect 925 1528 926 1532
rect 1262 1528 1265 1538
rect 1606 1532 1610 1536
rect 1822 1532 1825 1538
rect 1514 1528 1521 1531
rect 968 1503 970 1507
rect 974 1503 977 1507
rect 981 1503 984 1507
rect 650 1488 651 1492
rect 949 1488 950 1492
rect 102 1471 105 1481
rect 542 1478 553 1481
rect 886 1478 897 1481
rect 1234 1478 1241 1481
rect 94 1468 105 1471
rect 438 1468 465 1471
rect 1674 1468 1689 1471
rect 158 1458 166 1461
rect 458 1458 481 1461
rect 730 1458 746 1461
rect 838 1461 841 1468
rect 838 1458 849 1461
rect 970 1458 993 1461
rect 1022 1458 1042 1461
rect 1662 1458 1678 1461
rect 742 1457 746 1458
rect 1038 1457 1042 1458
rect 290 1438 293 1442
rect 456 1403 458 1407
rect 462 1403 465 1407
rect 469 1403 472 1407
rect 1480 1403 1482 1407
rect 1486 1403 1489 1407
rect 1493 1403 1496 1407
rect 508 1388 510 1392
rect 613 1388 614 1392
rect 780 1388 782 1392
rect 941 1388 942 1392
rect 1085 1388 1086 1392
rect 1149 1388 1150 1392
rect 1506 1368 1521 1371
rect 254 1348 262 1351
rect 598 1351 601 1361
rect 1630 1358 1638 1361
rect 582 1348 601 1351
rect 958 1348 966 1351
rect 1102 1348 1110 1351
rect 1166 1348 1174 1351
rect 1302 1348 1310 1351
rect 1342 1348 1353 1351
rect 1378 1348 1385 1351
rect 198 1341 201 1348
rect 198 1338 209 1341
rect 322 1338 329 1341
rect 438 1338 450 1341
rect 740 1338 742 1342
rect 850 1338 865 1341
rect 966 1341 969 1348
rect 1350 1342 1353 1348
rect 966 1338 993 1341
rect 1454 1341 1457 1348
rect 1842 1348 1857 1351
rect 1454 1338 1465 1341
rect 1486 1338 1505 1341
rect 1518 1338 1529 1341
rect 1674 1338 1681 1341
rect 1934 1338 1950 1341
rect 438 1332 441 1338
rect 710 1332 713 1338
rect 1502 1332 1505 1338
rect 242 1328 243 1332
rect 706 1328 713 1332
rect 878 1328 889 1331
rect 1506 1328 1513 1331
rect 1421 1318 1422 1322
rect 1450 1318 1451 1322
rect 1794 1318 1801 1321
rect 968 1303 970 1307
rect 974 1303 977 1307
rect 981 1303 984 1307
rect 458 1288 473 1291
rect 1690 1288 1692 1292
rect 594 1278 606 1281
rect 694 1278 713 1281
rect 718 1278 726 1281
rect 110 1272 114 1274
rect 141 1268 142 1272
rect 294 1262 297 1271
rect 682 1268 689 1271
rect 786 1268 793 1271
rect 870 1271 873 1281
rect 902 1278 914 1281
rect 1398 1278 1409 1281
rect 1450 1278 1465 1281
rect 1590 1278 1598 1282
rect 1630 1278 1641 1281
rect 1845 1278 1846 1282
rect 910 1277 914 1278
rect 1590 1272 1593 1278
rect 842 1268 849 1271
rect 854 1268 873 1271
rect 1354 1268 1361 1271
rect 1510 1268 1537 1271
rect 230 1258 238 1261
rect 318 1258 326 1261
rect 366 1258 374 1261
rect 590 1258 601 1261
rect 782 1258 798 1261
rect 850 1258 857 1261
rect 890 1258 897 1261
rect 1214 1258 1222 1261
rect 1446 1258 1454 1261
rect 1550 1258 1553 1268
rect 1630 1261 1633 1268
rect 1622 1258 1633 1261
rect 598 1252 601 1258
rect 326 1248 334 1251
rect 342 1248 353 1251
rect 446 1248 473 1251
rect 534 1248 545 1251
rect 618 1248 625 1251
rect 802 1248 806 1252
rect 814 1248 822 1251
rect 586 1238 587 1242
rect 778 1238 779 1242
rect 1590 1241 1594 1244
rect 1578 1238 1594 1241
rect 1746 1238 1749 1242
rect 365 1218 366 1222
rect 456 1203 458 1207
rect 462 1203 465 1207
rect 469 1203 472 1207
rect 1480 1203 1482 1207
rect 1486 1203 1489 1207
rect 1493 1203 1496 1207
rect 246 1188 257 1191
rect 1134 1188 1145 1191
rect 502 1171 505 1181
rect 502 1168 510 1171
rect 462 1158 478 1161
rect 550 1158 558 1161
rect 622 1158 630 1161
rect 594 1148 601 1151
rect 830 1151 833 1161
rect 830 1148 849 1151
rect 662 1138 673 1141
rect 790 1138 809 1141
rect 910 1141 913 1151
rect 1266 1148 1273 1151
rect 1382 1151 1385 1161
rect 1366 1148 1385 1151
rect 894 1138 913 1141
rect 1038 1138 1050 1141
rect 1246 1138 1254 1141
rect 1326 1138 1345 1141
rect 1406 1138 1417 1141
rect 670 1132 673 1138
rect 374 1128 385 1131
rect 558 1128 574 1131
rect 694 1131 698 1133
rect 690 1128 698 1131
rect 1438 1128 1454 1131
rect 1317 1118 1318 1122
rect 968 1103 970 1107
rect 974 1103 977 1107
rect 981 1103 984 1107
rect 1845 1088 1846 1092
rect 434 1078 446 1081
rect 450 1078 457 1081
rect 54 1068 65 1071
rect 222 1068 233 1071
rect 242 1068 249 1071
rect 350 1068 361 1071
rect 434 1068 465 1071
rect 734 1068 745 1071
rect 1534 1068 1545 1071
rect 1710 1068 1729 1071
rect 14 1058 33 1061
rect 46 1058 54 1061
rect 102 1058 110 1061
rect 182 1058 201 1061
rect 214 1058 222 1061
rect 310 1058 329 1061
rect 658 1058 665 1061
rect 726 1058 734 1061
rect 1134 1061 1137 1068
rect 1134 1058 1145 1061
rect 1406 1058 1414 1061
rect 1478 1058 1513 1061
rect 1562 1058 1569 1061
rect 1606 1058 1633 1061
rect 1710 1058 1718 1061
rect 1726 1058 1729 1068
rect 1862 1058 1870 1061
rect 30 1048 33 1058
rect 198 1048 201 1058
rect 326 1048 329 1058
rect 594 1048 601 1051
rect 1486 1048 1494 1051
rect 1510 1048 1513 1058
rect 378 1038 385 1041
rect 157 1018 158 1022
rect 562 1018 563 1022
rect 626 1018 627 1022
rect 1594 1018 1595 1022
rect 456 1003 458 1007
rect 462 1003 465 1007
rect 469 1003 472 1007
rect 1480 1003 1482 1007
rect 1486 1003 1489 1007
rect 1493 1003 1496 1007
rect 22 948 30 951
rect 46 948 54 951
rect 290 948 297 951
rect 318 948 329 951
rect 386 948 393 951
rect 482 948 508 951
rect 618 948 657 951
rect 766 948 774 951
rect 326 942 329 948
rect 54 938 65 941
rect 74 938 81 941
rect 130 938 138 941
rect 430 938 438 941
rect 454 938 462 941
rect 474 938 489 941
rect 578 938 585 941
rect 782 941 785 951
rect 854 941 857 951
rect 1166 951 1169 961
rect 1154 948 1169 951
rect 870 941 873 948
rect 694 938 705 941
rect 766 938 785 941
rect 838 938 857 941
rect 862 938 873 941
rect 1170 938 1177 941
rect 1230 938 1241 941
rect 1630 938 1642 941
rect 134 936 138 938
rect 390 931 393 938
rect 1430 932 1434 933
rect 382 928 393 931
rect 406 928 422 931
rect 1106 928 1107 932
rect 1314 928 1321 931
rect 108 918 110 922
rect 1284 918 1286 922
rect 1394 918 1396 922
rect 968 903 970 907
rect 974 903 977 907
rect 981 903 984 907
rect 18 888 19 892
rect 402 888 403 892
rect 516 888 518 892
rect 725 888 726 892
rect 1205 888 1206 892
rect 350 872 353 881
rect 378 878 385 882
rect 1242 878 1243 882
rect 1794 878 1801 881
rect 382 872 385 878
rect 1094 874 1098 878
rect 282 868 289 871
rect 310 868 329 871
rect 566 868 577 871
rect 742 871 746 874
rect 734 868 746 871
rect 1374 868 1382 871
rect 70 858 78 861
rect 110 858 118 861
rect 246 858 254 861
rect 302 861 305 868
rect 294 858 305 861
rect 558 858 566 861
rect 794 858 801 861
rect 1390 861 1393 868
rect 1390 858 1401 861
rect 1506 858 1513 861
rect 1598 858 1617 861
rect 1718 861 1721 868
rect 1710 858 1721 861
rect 1726 858 1742 861
rect 1806 861 1809 881
rect 1934 868 1942 871
rect 1806 858 1833 861
rect 354 848 361 851
rect 1598 848 1601 858
rect 1662 856 1666 858
rect 429 838 430 842
rect 602 838 609 841
rect 890 838 893 842
rect 1706 838 1707 842
rect 53 818 54 822
rect 1746 818 1747 822
rect 456 803 458 807
rect 462 803 465 807
rect 469 803 472 807
rect 1480 803 1482 807
rect 1486 803 1489 807
rect 1493 803 1496 807
rect 426 788 427 792
rect 510 761 513 768
rect 502 758 513 761
rect 554 758 558 762
rect 810 758 814 762
rect 822 758 830 761
rect 1694 758 1705 761
rect 1230 753 1234 758
rect 86 748 97 751
rect 94 742 97 748
rect 486 748 494 751
rect 1114 748 1121 751
rect 1574 748 1582 751
rect 1646 748 1654 751
rect 1706 748 1713 751
rect 1718 748 1753 751
rect 70 738 78 741
rect 190 738 202 741
rect 570 738 577 741
rect 886 741 889 748
rect 886 738 905 741
rect 1342 738 1350 741
rect 1386 738 1394 741
rect 1790 738 1817 741
rect 1822 738 1833 741
rect 450 728 470 731
rect 574 728 577 738
rect 1254 731 1257 738
rect 1630 732 1634 733
rect 1254 728 1265 731
rect 525 718 526 722
rect 1674 718 1675 722
rect 968 703 970 707
rect 974 703 977 707
rect 981 703 984 707
rect 478 688 486 691
rect 1002 688 1009 691
rect 566 678 577 681
rect 1110 678 1121 681
rect 1606 678 1614 682
rect 1690 678 1697 682
rect 1710 678 1718 681
rect 222 668 233 671
rect 366 668 377 671
rect 1038 668 1041 678
rect 1606 672 1609 678
rect 1694 672 1697 678
rect 1670 668 1681 671
rect 1934 668 1942 671
rect 214 658 222 661
rect 278 658 294 661
rect 358 658 366 661
rect 566 658 569 668
rect 758 658 766 661
rect 874 658 881 661
rect 1174 658 1190 661
rect 1510 658 1521 661
rect 1654 658 1673 661
rect 1710 658 1721 661
rect 1726 658 1734 661
rect 1770 658 1777 661
rect 534 651 537 658
rect 1654 656 1658 658
rect 510 648 521 651
rect 526 648 537 651
rect 1754 648 1758 652
rect 1867 638 1870 642
rect 478 618 486 621
rect 1781 618 1782 622
rect 456 603 458 607
rect 462 603 465 607
rect 469 603 472 607
rect 1480 603 1482 607
rect 1486 603 1489 607
rect 1493 603 1496 607
rect 262 548 278 551
rect 398 551 401 561
rect 486 558 505 561
rect 918 558 937 561
rect 1742 558 1753 561
rect 1646 552 1650 554
rect 378 548 385 551
rect 398 548 417 551
rect 450 548 473 551
rect 710 548 721 551
rect 894 548 913 551
rect 934 548 985 551
rect 1082 548 1090 551
rect 1514 548 1537 551
rect 1594 548 1601 551
rect 1754 548 1761 551
rect 710 542 713 548
rect 1086 546 1090 548
rect 170 538 185 541
rect 366 538 377 541
rect 438 538 465 541
rect 962 538 977 541
rect 1046 538 1089 541
rect 1194 538 1201 541
rect 1206 538 1214 541
rect 1334 538 1345 541
rect 1358 538 1385 541
rect 1414 538 1425 541
rect 1430 538 1457 541
rect 1474 538 1497 541
rect 1534 538 1545 541
rect 1786 538 1793 541
rect 86 528 94 531
rect 250 528 251 532
rect 778 528 779 532
rect 954 528 969 531
rect 1342 528 1345 538
rect 1470 528 1478 531
rect 1614 528 1617 538
rect 1910 532 1914 536
rect 1666 528 1681 531
rect 993 518 1014 521
rect 1562 518 1564 522
rect 968 503 970 507
rect 974 503 977 507
rect 981 503 984 507
rect 426 488 428 492
rect 1097 488 1118 491
rect 1149 488 1150 492
rect 1382 488 1390 491
rect 1558 488 1566 491
rect 854 478 865 481
rect 582 476 586 478
rect 878 472 881 481
rect 870 468 878 471
rect 998 468 1025 471
rect 1158 468 1177 471
rect 1286 468 1298 471
rect 134 458 142 461
rect 374 458 422 461
rect 662 458 673 461
rect 814 461 817 468
rect 1158 462 1161 468
rect 798 458 817 461
rect 822 458 841 461
rect 894 458 913 461
rect 1034 458 1041 461
rect 1526 461 1529 468
rect 1526 458 1537 461
rect 1706 458 1713 461
rect 1874 458 1881 461
rect 906 448 913 451
rect 1218 438 1221 442
rect 1602 438 1605 442
rect 456 403 458 407
rect 462 403 465 407
rect 469 403 472 407
rect 1480 403 1482 407
rect 1486 403 1489 407
rect 1493 403 1496 407
rect 434 388 435 392
rect 986 388 998 391
rect 786 368 793 371
rect 1867 368 1870 372
rect 146 348 161 351
rect 414 348 425 351
rect 462 348 481 351
rect 518 348 526 351
rect 566 348 574 351
rect 190 338 202 341
rect 326 332 329 342
rect 422 338 425 348
rect 462 341 465 348
rect 670 348 681 351
rect 702 351 705 361
rect 1142 353 1146 358
rect 698 348 705 351
rect 774 348 793 351
rect 830 348 846 351
rect 678 342 681 348
rect 1362 348 1369 351
rect 1606 348 1622 351
rect 1702 351 1706 353
rect 1694 348 1706 351
rect 454 338 465 341
rect 1050 338 1057 341
rect 1790 338 1802 341
rect 542 336 546 338
rect 1106 328 1113 331
rect 968 303 970 307
rect 974 303 977 307
rect 981 303 984 307
rect 1310 278 1321 281
rect 42 268 49 271
rect 142 268 145 278
rect 917 268 918 272
rect 1054 268 1057 278
rect 1622 274 1626 278
rect 1686 272 1690 274
rect 1450 268 1458 271
rect 710 258 718 261
rect 770 258 777 261
rect 1602 258 1609 261
rect 1662 258 1682 261
rect 1678 257 1682 258
rect 74 238 81 241
rect 1138 238 1141 242
rect 1411 238 1414 242
rect 742 228 745 238
rect 456 203 458 207
rect 462 203 465 207
rect 469 203 472 207
rect 1480 203 1482 207
rect 1486 203 1489 207
rect 1493 203 1496 207
rect 253 188 254 192
rect 1114 188 1115 192
rect 1518 188 1526 191
rect 370 168 373 172
rect 1499 168 1502 172
rect 786 158 793 161
rect 846 148 857 151
rect 1054 148 1081 151
rect 1118 148 1129 151
rect 782 138 790 141
rect 994 138 1001 141
rect 1042 138 1049 141
rect 1174 141 1177 148
rect 1190 141 1193 148
rect 1326 148 1345 151
rect 1142 138 1161 141
rect 1166 138 1177 141
rect 1182 138 1193 141
rect 1390 138 1393 148
rect 1622 148 1630 151
rect 1822 148 1830 151
rect 1586 138 1594 141
rect 1706 138 1713 141
rect 1726 138 1745 141
rect 1750 138 1769 141
rect 314 128 329 131
rect 334 128 342 131
rect 878 128 889 131
rect 998 128 1006 131
rect 1094 128 1105 131
rect 1214 131 1218 133
rect 1122 128 1129 131
rect 1190 128 1201 131
rect 1206 128 1218 131
rect 1230 132 1234 136
rect 1710 128 1713 138
rect 1058 118 1059 122
rect 968 103 970 107
rect 974 103 977 107
rect 981 103 984 107
rect 333 88 334 92
rect 1934 88 1942 91
rect 230 78 241 81
rect 246 78 270 81
rect 734 78 742 81
rect 1694 78 1705 81
rect 1710 78 1721 81
rect 1826 78 1833 81
rect 238 72 241 78
rect 734 77 738 78
rect 14 68 25 71
rect 62 68 86 71
rect 126 68 153 71
rect 302 68 310 71
rect 350 71 354 74
rect 342 68 354 71
rect 526 68 537 71
rect 1086 71 1090 74
rect 1078 68 1090 71
rect 1226 68 1233 71
rect 1374 71 1378 74
rect 1718 72 1721 78
rect 1374 68 1385 71
rect 126 61 129 68
rect 38 58 57 61
rect 110 58 129 61
rect 162 58 177 61
rect 458 58 473 61
rect 478 58 494 61
rect 538 58 545 61
rect 678 58 694 61
rect 750 58 761 61
rect 1234 58 1241 61
rect 1266 58 1273 61
rect 1674 58 1681 61
rect 546 48 550 52
rect 830 48 841 51
rect 1182 48 1185 58
rect 1502 38 1529 41
rect 456 3 458 7
rect 462 3 465 7
rect 469 3 472 7
rect 1480 3 1482 7
rect 1486 3 1489 7
rect 1493 3 1496 7
<< m2contact >>
rect 970 1703 974 1707
rect 977 1703 981 1707
rect 174 1688 178 1692
rect 222 1688 226 1692
rect 822 1688 826 1692
rect 870 1688 874 1692
rect 1062 1688 1066 1692
rect 1166 1688 1170 1692
rect 1206 1688 1210 1692
rect 1310 1688 1314 1692
rect 1350 1688 1354 1692
rect 1750 1688 1754 1692
rect 1854 1688 1858 1692
rect 1894 1688 1898 1692
rect 1918 1688 1922 1692
rect 70 1678 74 1682
rect 6 1668 10 1672
rect 30 1668 34 1672
rect 54 1668 58 1672
rect 62 1668 66 1672
rect 126 1678 130 1682
rect 198 1678 202 1682
rect 422 1678 426 1682
rect 622 1678 626 1682
rect 846 1678 850 1682
rect 902 1678 906 1682
rect 1022 1678 1026 1682
rect 1054 1679 1058 1683
rect 1454 1678 1458 1682
rect 1510 1678 1514 1682
rect 1862 1679 1866 1683
rect 1926 1678 1930 1682
rect 94 1668 98 1672
rect 118 1668 122 1672
rect 134 1668 138 1672
rect 142 1668 146 1672
rect 310 1668 314 1672
rect 406 1668 410 1672
rect 694 1668 698 1672
rect 806 1668 810 1672
rect 1150 1668 1154 1672
rect 1382 1668 1386 1672
rect 1606 1668 1610 1672
rect 1838 1668 1842 1672
rect 22 1658 26 1662
rect 78 1658 82 1662
rect 102 1658 106 1662
rect 150 1658 154 1662
rect 158 1658 162 1662
rect 182 1658 186 1662
rect 294 1659 298 1663
rect 390 1659 394 1663
rect 430 1658 434 1662
rect 438 1658 442 1662
rect 446 1658 450 1662
rect 470 1658 474 1662
rect 486 1658 490 1662
rect 494 1658 498 1662
rect 550 1658 554 1662
rect 574 1659 578 1663
rect 606 1658 610 1662
rect 622 1658 626 1662
rect 670 1658 674 1662
rect 790 1659 794 1663
rect 862 1658 866 1662
rect 886 1658 890 1662
rect 942 1658 946 1662
rect 974 1659 978 1663
rect 1014 1658 1018 1662
rect 1038 1658 1042 1662
rect 1046 1658 1050 1662
rect 1126 1658 1130 1662
rect 1182 1658 1186 1662
rect 1190 1658 1194 1662
rect 1246 1658 1250 1662
rect 1270 1658 1274 1662
rect 1326 1658 1330 1662
rect 1390 1658 1394 1662
rect 1454 1658 1458 1662
rect 1470 1658 1474 1662
rect 1494 1658 1498 1662
rect 1502 1658 1506 1662
rect 1526 1658 1530 1662
rect 1598 1658 1602 1662
rect 1670 1658 1674 1662
rect 1694 1658 1698 1662
rect 1734 1658 1738 1662
rect 1798 1658 1802 1662
rect 1814 1658 1818 1662
rect 1870 1658 1874 1662
rect 1878 1658 1882 1662
rect 1902 1658 1906 1662
rect 118 1648 122 1652
rect 1318 1638 1322 1642
rect 1742 1638 1746 1642
rect 1886 1638 1890 1642
rect 1910 1638 1914 1642
rect 230 1618 234 1622
rect 326 1618 330 1622
rect 510 1618 514 1622
rect 630 1618 634 1622
rect 726 1618 730 1622
rect 910 1618 914 1622
rect 1070 1618 1074 1622
rect 1214 1618 1218 1622
rect 1446 1618 1450 1622
rect 1542 1618 1546 1622
rect 1726 1618 1730 1622
rect 1758 1618 1762 1622
rect 1942 1618 1946 1622
rect 1926 1608 1930 1612
rect 458 1603 462 1607
rect 465 1603 469 1607
rect 1482 1603 1486 1607
rect 1489 1603 1493 1607
rect 126 1588 130 1592
rect 214 1588 218 1592
rect 262 1588 266 1592
rect 1070 1588 1074 1592
rect 1094 1588 1098 1592
rect 1118 1588 1122 1592
rect 1150 1588 1154 1592
rect 1270 1588 1274 1592
rect 1318 1588 1322 1592
rect 1622 1588 1626 1592
rect 1670 1588 1674 1592
rect 1814 1588 1818 1592
rect 1918 1578 1922 1582
rect 310 1568 314 1572
rect 822 1568 826 1572
rect 982 1568 986 1572
rect 1606 1568 1610 1572
rect 1790 1568 1794 1572
rect 1022 1558 1026 1562
rect 62 1548 66 1552
rect 102 1548 106 1552
rect 142 1548 146 1552
rect 158 1548 162 1552
rect 190 1548 194 1552
rect 206 1548 210 1552
rect 238 1548 242 1552
rect 254 1548 258 1552
rect 286 1548 290 1552
rect 358 1547 362 1551
rect 414 1547 418 1551
rect 550 1548 554 1552
rect 574 1548 578 1552
rect 670 1548 674 1552
rect 774 1547 778 1551
rect 870 1547 874 1551
rect 910 1548 914 1552
rect 942 1548 946 1552
rect 950 1548 954 1552
rect 1006 1548 1010 1552
rect 1014 1548 1018 1552
rect 1030 1548 1034 1552
rect 1078 1548 1082 1552
rect 1102 1548 1106 1552
rect 1110 1548 1114 1552
rect 1134 1548 1138 1552
rect 1222 1548 1226 1552
rect 1238 1548 1242 1552
rect 1254 1548 1258 1552
rect 1286 1548 1290 1552
rect 1294 1548 1298 1552
rect 1302 1548 1306 1552
rect 1326 1548 1330 1552
rect 1382 1548 1386 1552
rect 1406 1548 1410 1552
rect 1446 1548 1450 1552
rect 1454 1548 1458 1552
rect 1462 1548 1466 1552
rect 1478 1548 1482 1552
rect 1486 1548 1490 1552
rect 1502 1548 1506 1552
rect 1510 1548 1514 1552
rect 1566 1548 1570 1552
rect 1646 1548 1650 1552
rect 1662 1548 1666 1552
rect 150 1538 154 1542
rect 326 1538 330 1542
rect 374 1538 378 1542
rect 422 1538 426 1542
rect 598 1538 602 1542
rect 694 1538 698 1542
rect 886 1538 890 1542
rect 958 1538 962 1542
rect 1214 1538 1218 1542
rect 1254 1538 1258 1542
rect 1342 1538 1346 1542
rect 1542 1538 1546 1542
rect 1694 1548 1698 1552
rect 1718 1548 1722 1552
rect 1734 1548 1738 1552
rect 1742 1548 1746 1552
rect 1766 1548 1770 1552
rect 1774 1548 1778 1552
rect 1798 1548 1802 1552
rect 1806 1548 1810 1552
rect 1854 1547 1858 1551
rect 1926 1548 1930 1552
rect 1950 1538 1954 1542
rect 70 1528 74 1532
rect 510 1528 514 1532
rect 774 1528 778 1532
rect 926 1528 930 1532
rect 974 1528 978 1532
rect 1046 1528 1050 1532
rect 1174 1528 1178 1532
rect 1198 1528 1202 1532
rect 1278 1528 1282 1532
rect 1342 1528 1346 1532
rect 1510 1528 1514 1532
rect 1526 1528 1530 1532
rect 1606 1528 1610 1532
rect 1662 1528 1666 1532
rect 1822 1528 1826 1532
rect 6 1518 10 1522
rect 294 1518 298 1522
rect 478 1518 482 1522
rect 518 1518 522 1522
rect 614 1518 618 1522
rect 710 1518 714 1522
rect 806 1518 810 1522
rect 1350 1518 1354 1522
rect 1630 1518 1634 1522
rect 970 1503 974 1507
rect 977 1503 981 1507
rect 406 1488 410 1492
rect 614 1488 618 1492
rect 646 1488 650 1492
rect 686 1488 690 1492
rect 878 1488 882 1492
rect 950 1488 954 1492
rect 1014 1488 1018 1492
rect 1038 1488 1042 1492
rect 1134 1488 1138 1492
rect 1326 1488 1330 1492
rect 1478 1488 1482 1492
rect 1598 1488 1602 1492
rect 1622 1488 1626 1492
rect 86 1468 90 1472
rect 398 1478 402 1482
rect 534 1478 538 1482
rect 622 1478 626 1482
rect 710 1478 714 1482
rect 838 1478 842 1482
rect 1230 1478 1234 1482
rect 1246 1478 1250 1482
rect 1694 1478 1698 1482
rect 1718 1478 1722 1482
rect 1750 1478 1754 1482
rect 326 1468 330 1472
rect 374 1468 378 1472
rect 390 1468 394 1472
rect 414 1468 418 1472
rect 430 1468 434 1472
rect 510 1468 514 1472
rect 526 1468 530 1472
rect 574 1468 578 1472
rect 582 1468 586 1472
rect 606 1468 610 1472
rect 734 1468 738 1472
rect 774 1468 778 1472
rect 822 1468 826 1472
rect 838 1468 842 1472
rect 870 1468 874 1472
rect 918 1468 922 1472
rect 1214 1468 1218 1472
rect 1254 1468 1258 1472
rect 1318 1468 1322 1472
rect 1422 1468 1426 1472
rect 1518 1468 1522 1472
rect 1606 1468 1610 1472
rect 1670 1468 1674 1472
rect 1758 1468 1762 1472
rect 1830 1468 1834 1472
rect 62 1458 66 1462
rect 110 1458 114 1462
rect 118 1458 122 1462
rect 126 1458 130 1462
rect 134 1458 138 1462
rect 150 1458 154 1462
rect 166 1458 170 1462
rect 206 1458 210 1462
rect 238 1459 242 1463
rect 334 1459 338 1463
rect 382 1458 386 1462
rect 422 1458 426 1462
rect 454 1458 458 1462
rect 518 1458 522 1462
rect 566 1458 570 1462
rect 598 1458 602 1462
rect 630 1458 634 1462
rect 638 1458 642 1462
rect 662 1458 666 1462
rect 702 1458 706 1462
rect 726 1458 730 1462
rect 806 1459 810 1463
rect 854 1458 858 1462
rect 862 1458 866 1462
rect 910 1458 914 1462
rect 934 1458 938 1462
rect 966 1458 970 1462
rect 1070 1458 1074 1462
rect 1102 1459 1106 1463
rect 1198 1459 1202 1463
rect 1230 1458 1234 1462
rect 1358 1458 1362 1462
rect 1390 1459 1394 1463
rect 1542 1458 1546 1462
rect 1630 1458 1634 1462
rect 1638 1458 1642 1462
rect 1678 1458 1682 1462
rect 1702 1458 1706 1462
rect 1750 1459 1754 1463
rect 1846 1459 1850 1463
rect 1918 1458 1922 1462
rect 366 1448 370 1452
rect 550 1448 554 1452
rect 710 1448 714 1452
rect 894 1448 898 1452
rect 1622 1448 1626 1452
rect 1654 1448 1658 1452
rect 1710 1448 1714 1452
rect 6 1438 10 1442
rect 286 1438 290 1442
rect 1814 1428 1818 1432
rect 1910 1428 1914 1432
rect 174 1418 178 1422
rect 270 1418 274 1422
rect 438 1418 442 1422
rect 590 1418 594 1422
rect 742 1418 746 1422
rect 1134 1418 1138 1422
rect 1326 1418 1330 1422
rect 1614 1418 1618 1422
rect 458 1403 462 1407
rect 465 1403 469 1407
rect 1482 1403 1486 1407
rect 1489 1403 1493 1407
rect 510 1388 514 1392
rect 542 1388 546 1392
rect 614 1388 618 1392
rect 670 1388 674 1392
rect 782 1388 786 1392
rect 830 1388 834 1392
rect 942 1388 946 1392
rect 1038 1388 1042 1392
rect 1086 1388 1090 1392
rect 1150 1388 1154 1392
rect 1198 1388 1202 1392
rect 1238 1388 1242 1392
rect 1294 1388 1298 1392
rect 638 1378 642 1382
rect 6 1368 10 1372
rect 190 1368 194 1372
rect 446 1368 450 1372
rect 646 1368 650 1372
rect 678 1368 682 1372
rect 734 1368 738 1372
rect 1318 1368 1322 1372
rect 1502 1368 1506 1372
rect 1910 1368 1914 1372
rect 366 1358 370 1362
rect 430 1358 434 1362
rect 590 1358 594 1362
rect 62 1348 66 1352
rect 134 1348 138 1352
rect 198 1348 202 1352
rect 214 1348 218 1352
rect 222 1348 226 1352
rect 230 1348 234 1352
rect 262 1348 266 1352
rect 270 1348 274 1352
rect 294 1348 298 1352
rect 326 1348 330 1352
rect 350 1348 354 1352
rect 358 1348 362 1352
rect 382 1348 386 1352
rect 422 1348 426 1352
rect 446 1348 450 1352
rect 558 1348 562 1352
rect 574 1348 578 1352
rect 630 1358 634 1362
rect 662 1358 666 1362
rect 710 1358 714 1362
rect 718 1358 722 1362
rect 886 1358 890 1362
rect 1374 1358 1378 1362
rect 1414 1358 1418 1362
rect 1454 1358 1458 1362
rect 1462 1358 1466 1362
rect 1550 1358 1554 1362
rect 1638 1358 1642 1362
rect 614 1348 618 1352
rect 638 1348 642 1352
rect 670 1348 674 1352
rect 726 1348 730 1352
rect 806 1348 810 1352
rect 814 1348 818 1352
rect 838 1348 842 1352
rect 854 1348 858 1352
rect 902 1348 906 1352
rect 926 1348 930 1352
rect 966 1348 970 1352
rect 1006 1348 1010 1352
rect 1014 1348 1018 1352
rect 1046 1348 1050 1352
rect 1070 1348 1074 1352
rect 1110 1348 1114 1352
rect 1134 1348 1138 1352
rect 1174 1348 1178 1352
rect 1206 1348 1210 1352
rect 1230 1348 1234 1352
rect 1254 1348 1258 1352
rect 1262 1348 1266 1352
rect 1270 1348 1274 1352
rect 1278 1348 1282 1352
rect 1310 1348 1314 1352
rect 1358 1348 1362 1352
rect 1374 1348 1378 1352
rect 1454 1348 1458 1352
rect 1478 1348 1482 1352
rect 1534 1348 1538 1352
rect 1574 1348 1578 1352
rect 1614 1348 1618 1352
rect 1654 1348 1658 1352
rect 1694 1348 1698 1352
rect 70 1338 74 1342
rect 142 1338 146 1342
rect 318 1338 322 1342
rect 374 1338 378 1342
rect 390 1338 394 1342
rect 414 1338 418 1342
rect 478 1338 482 1342
rect 526 1338 530 1342
rect 566 1338 570 1342
rect 622 1338 626 1342
rect 694 1338 698 1342
rect 710 1338 714 1342
rect 742 1338 746 1342
rect 750 1338 754 1342
rect 798 1338 802 1342
rect 846 1338 850 1342
rect 910 1338 914 1342
rect 1334 1338 1338 1342
rect 1350 1338 1354 1342
rect 1374 1338 1378 1342
rect 1398 1338 1402 1342
rect 1430 1338 1434 1342
rect 1438 1338 1442 1342
rect 1726 1347 1730 1351
rect 1758 1348 1762 1352
rect 1830 1348 1834 1352
rect 1838 1348 1842 1352
rect 1894 1348 1898 1352
rect 1918 1348 1922 1352
rect 1558 1338 1562 1342
rect 1582 1338 1586 1342
rect 1606 1338 1610 1342
rect 1622 1338 1626 1342
rect 1646 1338 1650 1342
rect 1662 1338 1666 1342
rect 1670 1338 1674 1342
rect 1686 1338 1690 1342
rect 1950 1338 1954 1342
rect 198 1328 202 1332
rect 238 1328 242 1332
rect 278 1327 282 1331
rect 310 1328 314 1332
rect 398 1328 402 1332
rect 438 1328 442 1332
rect 1110 1328 1114 1332
rect 1318 1328 1322 1332
rect 1406 1328 1410 1332
rect 1502 1328 1506 1332
rect 1598 1328 1602 1332
rect 1670 1328 1674 1332
rect 1902 1327 1906 1331
rect 302 1318 306 1322
rect 406 1318 410 1322
rect 870 1318 874 1322
rect 1422 1318 1426 1322
rect 1446 1318 1450 1322
rect 1550 1318 1554 1322
rect 1566 1318 1570 1322
rect 1590 1318 1594 1322
rect 1790 1318 1794 1322
rect 970 1303 974 1307
rect 977 1303 981 1307
rect 286 1288 290 1292
rect 302 1288 306 1292
rect 454 1288 458 1292
rect 510 1288 514 1292
rect 654 1288 658 1292
rect 718 1288 722 1292
rect 822 1288 826 1292
rect 878 1288 882 1292
rect 1030 1288 1034 1292
rect 1102 1288 1106 1292
rect 1342 1288 1346 1292
rect 1470 1288 1474 1292
rect 1686 1288 1690 1292
rect 334 1278 338 1282
rect 382 1278 386 1282
rect 438 1278 442 1282
rect 518 1278 522 1282
rect 526 1278 530 1282
rect 574 1278 578 1282
rect 590 1278 594 1282
rect 726 1278 730 1282
rect 766 1278 770 1282
rect 86 1268 90 1272
rect 110 1268 114 1272
rect 142 1268 146 1272
rect 182 1268 186 1272
rect 62 1258 66 1262
rect 166 1259 170 1263
rect 310 1268 314 1272
rect 374 1268 378 1272
rect 494 1268 498 1272
rect 614 1268 618 1272
rect 638 1268 642 1272
rect 678 1268 682 1272
rect 718 1268 722 1272
rect 782 1268 786 1272
rect 838 1268 842 1272
rect 1174 1278 1178 1282
rect 1198 1278 1202 1282
rect 1518 1278 1522 1282
rect 1550 1278 1554 1282
rect 1846 1278 1850 1282
rect 1870 1278 1874 1282
rect 1886 1278 1890 1282
rect 1934 1278 1938 1282
rect 990 1268 994 1272
rect 1086 1268 1090 1272
rect 1222 1268 1226 1272
rect 1350 1268 1354 1272
rect 1366 1268 1370 1272
rect 1374 1268 1378 1272
rect 1422 1268 1426 1272
rect 1438 1268 1442 1272
rect 1550 1268 1554 1272
rect 1590 1268 1594 1272
rect 1606 1268 1610 1272
rect 1630 1268 1634 1272
rect 1662 1268 1666 1272
rect 1670 1268 1674 1272
rect 1718 1268 1722 1272
rect 238 1258 242 1262
rect 254 1258 258 1262
rect 294 1258 298 1262
rect 326 1258 330 1262
rect 374 1258 378 1262
rect 398 1258 402 1262
rect 422 1258 426 1262
rect 486 1258 490 1262
rect 502 1258 506 1262
rect 550 1258 554 1262
rect 662 1258 666 1262
rect 678 1258 682 1262
rect 726 1258 730 1262
rect 798 1258 802 1262
rect 846 1258 850 1262
rect 886 1258 890 1262
rect 966 1258 970 1262
rect 1118 1258 1122 1262
rect 1126 1258 1130 1262
rect 1134 1258 1138 1262
rect 1158 1258 1162 1262
rect 1222 1258 1226 1262
rect 1294 1258 1298 1262
rect 1326 1258 1330 1262
rect 1382 1258 1386 1262
rect 1414 1258 1418 1262
rect 1430 1258 1434 1262
rect 1454 1258 1458 1262
rect 1478 1258 1482 1262
rect 1502 1258 1506 1262
rect 1526 1258 1530 1262
rect 1574 1258 1578 1262
rect 1614 1258 1618 1262
rect 1654 1258 1658 1262
rect 1758 1258 1762 1262
rect 1782 1258 1786 1262
rect 1830 1258 1834 1262
rect 1862 1258 1866 1262
rect 1894 1258 1898 1262
rect 1902 1258 1906 1262
rect 1910 1258 1914 1262
rect 1950 1258 1954 1262
rect 334 1248 338 1252
rect 430 1248 434 1252
rect 598 1248 602 1252
rect 614 1248 618 1252
rect 630 1248 634 1252
rect 670 1248 674 1252
rect 798 1248 802 1252
rect 822 1248 826 1252
rect 1398 1248 1402 1252
rect 1454 1248 1458 1252
rect 1558 1248 1562 1252
rect 1582 1248 1586 1252
rect 1638 1248 1642 1252
rect 6 1238 10 1242
rect 398 1238 402 1242
rect 414 1238 418 1242
rect 558 1238 562 1242
rect 582 1238 586 1242
rect 654 1238 658 1242
rect 774 1238 778 1242
rect 1566 1238 1570 1242
rect 1574 1238 1578 1242
rect 1742 1238 1746 1242
rect 1926 1238 1930 1242
rect 422 1228 426 1232
rect 910 1228 914 1232
rect 102 1218 106 1222
rect 286 1218 290 1222
rect 366 1218 370 1222
rect 502 1218 506 1222
rect 550 1218 554 1222
rect 1150 1218 1154 1222
rect 1278 1218 1282 1222
rect 1310 1218 1314 1222
rect 1502 1218 1506 1222
rect 1726 1218 1730 1222
rect 1950 1218 1954 1222
rect 458 1203 462 1207
rect 465 1203 469 1207
rect 1482 1203 1486 1207
rect 1489 1203 1493 1207
rect 6 1188 10 1192
rect 438 1188 442 1192
rect 694 1188 698 1192
rect 1430 1188 1434 1192
rect 430 1168 434 1172
rect 446 1168 450 1172
rect 494 1168 498 1172
rect 518 1178 522 1182
rect 510 1168 514 1172
rect 526 1168 530 1172
rect 1142 1168 1146 1172
rect 1686 1168 1690 1172
rect 1878 1168 1882 1172
rect 374 1158 378 1162
rect 478 1158 482 1162
rect 510 1158 514 1162
rect 542 1158 546 1162
rect 558 1158 562 1162
rect 566 1158 570 1162
rect 590 1158 594 1162
rect 630 1158 634 1162
rect 62 1148 66 1152
rect 118 1148 122 1152
rect 190 1148 194 1152
rect 286 1148 290 1152
rect 318 1147 322 1151
rect 358 1148 362 1152
rect 406 1148 410 1152
rect 430 1148 434 1152
rect 454 1148 458 1152
rect 502 1148 506 1152
rect 534 1148 538 1152
rect 590 1148 594 1152
rect 606 1148 610 1152
rect 654 1148 658 1152
rect 686 1148 690 1152
rect 758 1147 762 1151
rect 814 1148 818 1152
rect 838 1158 842 1162
rect 1278 1158 1282 1162
rect 1310 1158 1314 1162
rect 1374 1158 1378 1162
rect 862 1148 866 1152
rect 870 1148 874 1152
rect 894 1148 898 1152
rect 70 1138 74 1142
rect 126 1138 130 1142
rect 134 1140 138 1144
rect 350 1138 354 1142
rect 398 1138 402 1142
rect 582 1138 586 1142
rect 614 1138 618 1142
rect 774 1138 778 1142
rect 854 1138 858 1142
rect 1014 1147 1018 1151
rect 1078 1148 1082 1152
rect 1102 1148 1106 1152
rect 1174 1148 1178 1152
rect 1206 1147 1210 1151
rect 1254 1148 1258 1152
rect 1262 1148 1266 1152
rect 1294 1148 1298 1152
rect 1302 1148 1306 1152
rect 1350 1148 1354 1152
rect 1798 1158 1802 1162
rect 1830 1158 1834 1162
rect 1398 1148 1402 1152
rect 1526 1147 1530 1151
rect 1566 1148 1570 1152
rect 1654 1147 1658 1151
rect 1750 1147 1754 1151
rect 1790 1148 1794 1152
rect 1822 1148 1826 1152
rect 1838 1148 1842 1152
rect 1846 1148 1850 1152
rect 1862 1148 1866 1152
rect 1886 1148 1890 1152
rect 1902 1148 1906 1152
rect 1918 1148 1922 1152
rect 982 1138 986 1142
rect 1254 1138 1258 1142
rect 1358 1138 1362 1142
rect 1542 1138 1546 1142
rect 1558 1138 1562 1142
rect 1670 1138 1674 1142
rect 1766 1138 1770 1142
rect 1854 1138 1858 1142
rect 1894 1138 1898 1142
rect 102 1128 106 1132
rect 182 1128 186 1132
rect 390 1128 394 1132
rect 414 1128 418 1132
rect 574 1128 578 1132
rect 630 1128 634 1132
rect 670 1128 674 1132
rect 686 1128 690 1132
rect 798 1128 802 1132
rect 926 1128 930 1132
rect 1238 1128 1242 1132
rect 1334 1128 1338 1132
rect 1422 1128 1426 1132
rect 1454 1128 1458 1132
rect 1910 1128 1914 1132
rect 110 1118 114 1122
rect 150 1118 154 1122
rect 254 1118 258 1122
rect 638 1118 642 1122
rect 678 1118 682 1122
rect 918 1118 922 1122
rect 950 1118 954 1122
rect 1318 1118 1322 1122
rect 1462 1118 1466 1122
rect 1582 1118 1586 1122
rect 1590 1118 1594 1122
rect 970 1103 974 1107
rect 977 1103 981 1107
rect 1918 1098 1922 1102
rect 462 1088 466 1092
rect 702 1088 706 1092
rect 766 1088 770 1092
rect 830 1088 834 1092
rect 942 1088 946 1092
rect 1038 1088 1042 1092
rect 1166 1088 1170 1092
rect 1366 1088 1370 1092
rect 1462 1088 1466 1092
rect 1646 1088 1650 1092
rect 1734 1088 1738 1092
rect 1806 1088 1810 1092
rect 1846 1088 1850 1092
rect 1894 1088 1898 1092
rect 70 1078 74 1082
rect 110 1078 114 1082
rect 238 1078 242 1082
rect 366 1078 370 1082
rect 430 1078 434 1082
rect 446 1078 450 1082
rect 654 1078 658 1082
rect 750 1078 754 1082
rect 1134 1078 1138 1082
rect 1550 1078 1554 1082
rect 1558 1078 1562 1082
rect 1622 1078 1626 1082
rect 1742 1078 1746 1082
rect 1918 1078 1922 1082
rect 6 1068 10 1072
rect 78 1068 82 1072
rect 86 1066 90 1070
rect 134 1068 138 1072
rect 166 1068 170 1072
rect 174 1068 178 1072
rect 238 1068 242 1072
rect 294 1068 298 1072
rect 302 1068 306 1072
rect 374 1068 378 1072
rect 430 1068 434 1072
rect 590 1068 594 1072
rect 614 1068 618 1072
rect 646 1068 650 1072
rect 678 1068 682 1072
rect 686 1066 690 1070
rect 822 1068 826 1072
rect 910 1068 914 1072
rect 990 1068 994 1072
rect 1022 1068 1026 1072
rect 1134 1068 1138 1072
rect 1222 1068 1226 1072
rect 1286 1068 1290 1072
rect 1382 1068 1386 1072
rect 1470 1068 1474 1072
rect 1582 1068 1586 1072
rect 1614 1068 1618 1072
rect 1670 1068 1674 1072
rect 1750 1068 1754 1072
rect 54 1058 58 1062
rect 110 1058 114 1062
rect 126 1058 130 1062
rect 142 1058 146 1062
rect 158 1058 162 1062
rect 222 1058 226 1062
rect 342 1058 346 1062
rect 406 1058 410 1062
rect 470 1058 474 1062
rect 534 1058 538 1062
rect 542 1058 546 1062
rect 550 1058 554 1062
rect 574 1058 578 1062
rect 622 1058 626 1062
rect 638 1058 642 1062
rect 654 1058 658 1062
rect 670 1058 674 1062
rect 734 1058 738 1062
rect 894 1059 898 1063
rect 998 1058 1002 1062
rect 1070 1058 1074 1062
rect 1102 1059 1106 1063
rect 1150 1058 1154 1062
rect 1230 1058 1234 1062
rect 1238 1058 1242 1062
rect 1262 1058 1266 1062
rect 1310 1058 1314 1062
rect 1414 1058 1418 1062
rect 1526 1058 1530 1062
rect 1558 1058 1562 1062
rect 1574 1058 1578 1062
rect 1590 1058 1594 1062
rect 1638 1058 1642 1062
rect 1662 1058 1666 1062
rect 1678 1058 1682 1062
rect 1686 1058 1690 1062
rect 1718 1058 1722 1062
rect 1830 1058 1834 1062
rect 1870 1058 1874 1062
rect 1902 1058 1906 1062
rect 22 1048 26 1052
rect 190 1048 194 1052
rect 318 1048 322 1052
rect 390 1048 394 1052
rect 398 1048 402 1052
rect 590 1048 594 1052
rect 606 1048 610 1052
rect 710 1048 714 1052
rect 1494 1048 1498 1052
rect 126 1038 130 1042
rect 374 1038 378 1042
rect 414 1038 418 1042
rect 406 1028 410 1032
rect 158 1018 162 1022
rect 270 1018 274 1022
rect 518 1018 522 1022
rect 558 1018 562 1022
rect 622 1018 626 1022
rect 1254 1018 1258 1022
rect 1590 1018 1594 1022
rect 1806 1018 1810 1022
rect 458 1003 462 1007
rect 465 1003 469 1007
rect 1482 1003 1486 1007
rect 1489 1003 1493 1007
rect 134 988 138 992
rect 1046 988 1050 992
rect 1430 988 1434 992
rect 1542 988 1546 992
rect 878 978 882 982
rect 1190 978 1194 982
rect 1726 968 1730 972
rect 30 958 34 962
rect 350 958 354 962
rect 382 958 386 962
rect 414 958 418 962
rect 542 958 546 962
rect 726 958 730 962
rect 1134 958 1138 962
rect 30 948 34 952
rect 54 948 58 952
rect 166 948 170 952
rect 198 947 202 951
rect 262 948 266 952
rect 286 948 290 952
rect 334 948 338 952
rect 366 948 370 952
rect 382 948 386 952
rect 398 948 402 952
rect 462 948 466 952
rect 478 948 482 952
rect 590 948 594 952
rect 614 948 618 952
rect 710 948 714 952
rect 734 948 738 952
rect 742 948 746 952
rect 774 948 778 952
rect 6 938 10 942
rect 70 938 74 942
rect 126 938 130 942
rect 182 938 186 942
rect 254 938 258 942
rect 270 938 274 942
rect 310 938 314 942
rect 326 938 330 942
rect 342 938 346 942
rect 358 938 362 942
rect 390 938 394 942
rect 438 938 442 942
rect 462 938 466 942
rect 470 938 474 942
rect 534 938 538 942
rect 558 938 562 942
rect 574 938 578 942
rect 630 938 634 942
rect 678 938 682 942
rect 806 948 810 952
rect 814 948 818 952
rect 838 948 842 952
rect 870 948 874 952
rect 910 948 914 952
rect 934 948 938 952
rect 1078 948 1082 952
rect 1086 948 1090 952
rect 1094 948 1098 952
rect 1118 948 1122 952
rect 1150 948 1154 952
rect 1206 958 1210 962
rect 1222 948 1226 952
rect 1334 948 1338 952
rect 1494 947 1498 951
rect 1598 948 1602 952
rect 1662 947 1666 951
rect 1694 948 1698 952
rect 1766 948 1770 952
rect 1790 948 1794 952
rect 1854 947 1858 951
rect 1926 948 1930 952
rect 990 938 994 942
rect 1158 938 1162 942
rect 1166 938 1170 942
rect 1182 938 1186 942
rect 1254 938 1258 942
rect 1302 938 1306 942
rect 1334 938 1338 942
rect 1374 938 1378 942
rect 1422 938 1426 942
rect 1510 938 1514 942
rect 1838 938 1842 942
rect 1942 938 1946 942
rect 70 928 74 932
rect 270 928 274 932
rect 294 928 298 932
rect 438 928 442 932
rect 582 928 586 932
rect 686 928 690 932
rect 798 928 802 932
rect 870 928 874 932
rect 1062 928 1066 932
rect 1102 928 1106 932
rect 1198 928 1202 932
rect 1246 928 1250 932
rect 1310 928 1314 932
rect 1430 928 1434 932
rect 110 918 114 922
rect 446 918 450 922
rect 542 918 546 922
rect 582 918 586 922
rect 790 918 794 922
rect 878 918 882 922
rect 1046 918 1050 922
rect 1070 918 1074 922
rect 1286 918 1290 922
rect 1326 918 1330 922
rect 1390 918 1394 922
rect 1734 918 1738 922
rect 1918 918 1922 922
rect 1550 908 1554 912
rect 970 903 974 907
rect 977 903 981 907
rect 1926 898 1930 902
rect 14 888 18 892
rect 126 888 130 892
rect 230 888 234 892
rect 270 888 274 892
rect 342 888 346 892
rect 398 888 402 892
rect 454 888 458 892
rect 518 888 522 892
rect 622 888 626 892
rect 726 888 730 892
rect 742 888 746 892
rect 846 888 850 892
rect 870 888 874 892
rect 1206 888 1210 892
rect 1270 888 1274 892
rect 1454 888 1458 892
rect 1598 888 1602 892
rect 318 878 322 882
rect 446 878 450 882
rect 582 878 586 882
rect 1094 878 1098 882
rect 1174 878 1178 882
rect 1238 878 1242 882
rect 1366 878 1370 882
rect 1694 878 1698 882
rect 1766 878 1770 882
rect 1790 878 1794 882
rect 6 868 10 872
rect 182 868 186 872
rect 278 868 282 872
rect 302 868 306 872
rect 350 868 354 872
rect 366 868 370 872
rect 382 868 386 872
rect 390 868 394 872
rect 438 868 442 872
rect 486 868 490 872
rect 534 868 538 872
rect 702 868 706 872
rect 822 868 826 872
rect 950 868 954 872
rect 1062 868 1066 872
rect 1214 868 1218 872
rect 1334 868 1338 872
rect 1350 868 1354 872
rect 1382 868 1386 872
rect 1390 868 1394 872
rect 1510 868 1514 872
rect 1574 868 1578 872
rect 1622 868 1626 872
rect 1718 868 1722 872
rect 1734 868 1738 872
rect 38 858 42 862
rect 62 858 66 862
rect 78 858 82 862
rect 86 858 90 862
rect 118 858 122 862
rect 190 859 194 863
rect 254 858 258 862
rect 430 858 434 862
rect 462 858 466 862
rect 566 858 570 862
rect 598 858 602 862
rect 686 859 690 863
rect 790 858 794 862
rect 862 858 866 862
rect 934 859 938 863
rect 1046 859 1050 863
rect 1110 858 1114 862
rect 1134 858 1138 862
rect 1190 858 1194 862
rect 1222 858 1226 862
rect 1230 858 1234 862
rect 1254 858 1258 862
rect 1326 858 1330 862
rect 1382 858 1386 862
rect 1422 858 1426 862
rect 1430 858 1434 862
rect 1502 858 1506 862
rect 1550 858 1554 862
rect 1582 858 1586 862
rect 1646 858 1650 862
rect 1662 858 1666 862
rect 1678 858 1682 862
rect 1742 858 1746 862
rect 1782 858 1786 862
rect 1790 858 1794 862
rect 1902 879 1906 883
rect 1814 868 1818 872
rect 1862 868 1866 872
rect 1942 868 1946 872
rect 1886 858 1890 862
rect 1894 858 1898 862
rect 1918 858 1922 862
rect 22 848 26 852
rect 342 848 346 852
rect 350 848 354 852
rect 382 848 386 852
rect 406 848 410 852
rect 414 848 418 852
rect 542 848 546 852
rect 590 848 594 852
rect 718 848 722 852
rect 1198 848 1202 852
rect 1406 848 1410 852
rect 1606 848 1610 852
rect 1654 848 1658 852
rect 1758 848 1762 852
rect 430 838 434 842
rect 598 838 602 842
rect 886 838 890 842
rect 1638 838 1642 842
rect 1678 838 1682 842
rect 1702 838 1706 842
rect 1878 838 1882 842
rect 54 818 58 822
rect 102 818 106 822
rect 614 818 618 822
rect 982 818 986 822
rect 1078 818 1082 822
rect 1190 818 1194 822
rect 1646 818 1650 822
rect 1670 818 1674 822
rect 1742 818 1746 822
rect 1782 818 1786 822
rect 458 803 462 807
rect 465 803 469 807
rect 1482 803 1486 807
rect 1489 803 1493 807
rect 102 788 106 792
rect 286 788 290 792
rect 318 788 322 792
rect 422 788 426 792
rect 598 788 602 792
rect 1006 788 1010 792
rect 1030 788 1034 792
rect 1150 788 1154 792
rect 1374 788 1378 792
rect 1534 788 1538 792
rect 1630 788 1634 792
rect 654 778 658 782
rect 510 768 514 772
rect 646 768 650 772
rect 454 758 458 762
rect 518 758 522 762
rect 542 758 546 762
rect 558 758 562 762
rect 662 758 666 762
rect 806 758 810 762
rect 830 758 834 762
rect 862 758 866 762
rect 1230 758 1234 762
rect 1678 758 1682 762
rect 1806 758 1810 762
rect 78 748 82 752
rect 158 748 162 752
rect 230 748 234 752
rect 310 748 314 752
rect 382 747 386 751
rect 430 748 434 752
rect 478 748 482 752
rect 494 748 498 752
rect 558 748 562 752
rect 606 748 610 752
rect 654 748 658 752
rect 702 748 706 752
rect 734 747 738 751
rect 766 748 770 752
rect 806 748 810 752
rect 846 748 850 752
rect 878 748 882 752
rect 886 748 890 752
rect 918 748 922 752
rect 934 748 938 752
rect 958 748 962 752
rect 966 748 970 752
rect 990 748 994 752
rect 1094 748 1098 752
rect 1110 748 1114 752
rect 1190 748 1194 752
rect 1214 748 1218 752
rect 1254 748 1258 752
rect 1422 748 1426 752
rect 1502 748 1506 752
rect 1582 748 1586 752
rect 1638 748 1642 752
rect 1654 748 1658 752
rect 1702 748 1706 752
rect 1798 748 1802 752
rect 6 738 10 742
rect 78 738 82 742
rect 94 738 98 742
rect 150 738 154 742
rect 374 738 378 742
rect 438 738 442 742
rect 534 738 538 742
rect 566 738 570 742
rect 582 738 586 742
rect 614 738 618 742
rect 774 738 778 742
rect 798 738 802 742
rect 854 738 858 742
rect 1870 747 1874 751
rect 1054 738 1058 742
rect 1254 738 1258 742
rect 1278 738 1282 742
rect 1350 738 1354 742
rect 1382 738 1386 742
rect 1550 738 1554 742
rect 1662 738 1666 742
rect 1726 738 1730 742
rect 1854 738 1858 742
rect 94 728 98 732
rect 294 728 298 732
rect 414 728 418 732
rect 470 728 474 732
rect 494 728 498 732
rect 510 728 514 732
rect 630 728 634 732
rect 782 728 786 732
rect 790 728 794 732
rect 830 728 834 732
rect 1270 728 1274 732
rect 1526 728 1530 732
rect 1630 728 1634 732
rect 1654 728 1658 732
rect 1686 728 1690 732
rect 1734 728 1738 732
rect 1766 728 1770 732
rect 1774 728 1778 732
rect 1838 728 1842 732
rect 102 718 106 722
rect 302 718 306 722
rect 318 718 322 722
rect 526 718 530 722
rect 598 718 602 722
rect 622 718 626 722
rect 670 718 674 722
rect 862 718 866 722
rect 942 718 946 722
rect 1246 718 1250 722
rect 1478 718 1482 722
rect 1670 718 1674 722
rect 1758 718 1762 722
rect 1782 718 1786 722
rect 1934 718 1938 722
rect 22 708 26 712
rect 970 703 974 707
rect 977 703 981 707
rect 102 688 106 692
rect 334 688 338 692
rect 486 688 490 692
rect 630 688 634 692
rect 774 688 778 692
rect 982 688 986 692
rect 998 688 1002 692
rect 1398 688 1402 692
rect 1462 688 1466 692
rect 1638 688 1642 692
rect 1886 688 1890 692
rect 238 678 242 682
rect 382 678 386 682
rect 502 678 506 682
rect 622 678 626 682
rect 838 678 842 682
rect 870 678 874 682
rect 1038 678 1042 682
rect 1070 678 1074 682
rect 1166 678 1170 682
rect 1334 678 1338 682
rect 1718 678 1722 682
rect 1734 678 1738 682
rect 1790 678 1794 682
rect 30 668 34 672
rect 94 668 98 672
rect 182 668 186 672
rect 270 668 274 672
rect 398 668 402 672
rect 534 668 538 672
rect 550 668 554 672
rect 566 668 570 672
rect 598 668 602 672
rect 710 668 714 672
rect 934 668 938 672
rect 1238 668 1242 672
rect 1406 668 1410 672
rect 1542 668 1546 672
rect 1598 668 1602 672
rect 1606 668 1610 672
rect 1622 668 1626 672
rect 1662 668 1666 672
rect 1694 668 1698 672
rect 1702 668 1706 672
rect 1766 668 1770 672
rect 1806 668 1810 672
rect 1942 668 1946 672
rect 22 658 26 662
rect 166 659 170 663
rect 222 658 226 662
rect 294 658 298 662
rect 366 658 370 662
rect 422 658 426 662
rect 534 658 538 662
rect 542 658 546 662
rect 590 658 594 662
rect 606 658 610 662
rect 694 659 698 663
rect 726 658 730 662
rect 734 658 738 662
rect 766 658 770 662
rect 838 659 842 663
rect 870 658 874 662
rect 886 658 890 662
rect 918 659 922 663
rect 1070 659 1074 663
rect 1134 658 1138 662
rect 1190 658 1194 662
rect 1342 658 1346 662
rect 1534 658 1538 662
rect 1550 658 1554 662
rect 1590 658 1594 662
rect 1646 658 1650 662
rect 1734 658 1738 662
rect 1758 658 1762 662
rect 1766 658 1770 662
rect 1822 659 1826 663
rect 1894 658 1898 662
rect 1918 658 1922 662
rect 198 648 202 652
rect 342 648 346 652
rect 574 648 578 652
rect 1606 648 1610 652
rect 1694 648 1698 652
rect 1742 648 1746 652
rect 1758 648 1762 652
rect 6 638 10 642
rect 1230 638 1234 642
rect 1502 638 1506 642
rect 1638 638 1642 642
rect 1870 638 1874 642
rect 1902 638 1906 642
rect 1910 638 1914 642
rect 86 618 90 622
rect 486 618 490 622
rect 606 618 610 622
rect 750 618 754 622
rect 1294 618 1298 622
rect 1398 618 1402 622
rect 1670 618 1674 622
rect 1782 618 1786 622
rect 458 603 462 607
rect 465 603 469 607
rect 1482 603 1486 607
rect 1489 603 1493 607
rect 1918 598 1922 602
rect 158 588 162 592
rect 182 588 186 592
rect 286 588 290 592
rect 1110 588 1114 592
rect 1470 588 1474 592
rect 1622 588 1626 592
rect 1926 588 1930 592
rect 1934 588 1938 592
rect 1710 578 1714 582
rect 126 568 130 572
rect 518 568 522 572
rect 614 568 618 572
rect 1630 568 1634 572
rect 1718 568 1722 572
rect 166 558 170 562
rect 294 558 298 562
rect 94 548 98 552
rect 102 548 106 552
rect 110 548 114 552
rect 134 548 138 552
rect 198 548 202 552
rect 222 548 226 552
rect 230 548 234 552
rect 238 548 242 552
rect 278 548 282 552
rect 374 548 378 552
rect 406 558 410 562
rect 510 558 514 562
rect 830 558 834 562
rect 1158 558 1162 562
rect 1438 558 1442 562
rect 1494 558 1498 562
rect 1606 558 1610 562
rect 1670 558 1674 562
rect 1702 558 1706 562
rect 1806 558 1810 562
rect 446 548 450 552
rect 582 547 586 551
rect 646 548 650 552
rect 678 547 682 551
rect 726 548 730 552
rect 750 548 754 552
rect 758 548 762 552
rect 766 548 770 552
rect 790 548 794 552
rect 806 548 810 552
rect 838 548 842 552
rect 870 548 874 552
rect 886 548 890 552
rect 1038 548 1042 552
rect 1054 548 1058 552
rect 1062 548 1066 552
rect 1078 548 1082 552
rect 1094 548 1098 552
rect 1118 548 1122 552
rect 1134 548 1138 552
rect 1190 548 1194 552
rect 1222 548 1226 552
rect 1302 548 1306 552
rect 1366 548 1370 552
rect 1446 548 1450 552
rect 1510 548 1514 552
rect 1590 548 1594 552
rect 1638 548 1642 552
rect 1646 548 1650 552
rect 1694 548 1698 552
rect 1710 548 1714 552
rect 1750 548 1754 552
rect 1766 548 1770 552
rect 1798 548 1802 552
rect 1822 548 1826 552
rect 1862 547 1866 551
rect 6 538 10 542
rect 150 538 154 542
rect 166 538 170 542
rect 278 538 282 542
rect 302 538 306 542
rect 350 538 354 542
rect 422 538 426 542
rect 494 538 498 542
rect 574 538 578 542
rect 710 538 714 542
rect 862 538 866 542
rect 902 538 906 542
rect 958 538 962 542
rect 1030 538 1034 542
rect 1126 538 1130 542
rect 1142 538 1146 542
rect 1174 538 1178 542
rect 1190 538 1194 542
rect 1214 538 1218 542
rect 1278 538 1282 542
rect 1294 538 1298 542
rect 1390 538 1394 542
rect 1470 538 1474 542
rect 1518 538 1522 542
rect 1526 538 1530 542
rect 1614 538 1618 542
rect 1654 538 1658 542
rect 1774 538 1778 542
rect 1782 538 1786 542
rect 1830 538 1834 542
rect 1870 538 1874 542
rect 78 528 82 532
rect 94 528 98 532
rect 206 528 210 532
rect 246 528 250 532
rect 358 528 362 532
rect 430 528 434 532
rect 710 528 714 532
rect 734 528 738 532
rect 774 528 778 532
rect 846 528 850 532
rect 878 528 882 532
rect 926 528 930 532
rect 950 528 954 532
rect 1078 528 1082 532
rect 1182 528 1186 532
rect 1214 528 1218 532
rect 1374 528 1378 532
rect 1406 528 1410 532
rect 1478 528 1482 532
rect 1734 528 1738 532
rect 1782 528 1786 532
rect 1910 528 1914 532
rect 1942 528 1946 532
rect 62 518 66 522
rect 214 518 218 522
rect 326 518 330 522
rect 742 518 746 522
rect 854 518 858 522
rect 974 518 978 522
rect 1014 518 1018 522
rect 1246 518 1250 522
rect 1350 518 1354 522
rect 1558 518 1562 522
rect 1686 518 1690 522
rect 1806 518 1810 522
rect 22 508 26 512
rect 1918 508 1922 512
rect 970 503 974 507
rect 977 503 981 507
rect 30 488 34 492
rect 238 488 242 492
rect 334 488 338 492
rect 382 488 386 492
rect 422 488 426 492
rect 478 488 482 492
rect 686 488 690 492
rect 782 488 786 492
rect 862 488 866 492
rect 886 488 890 492
rect 934 488 938 492
rect 998 488 1002 492
rect 1118 488 1122 492
rect 1150 488 1154 492
rect 1182 488 1186 492
rect 1198 488 1202 492
rect 1390 488 1394 492
rect 1566 488 1570 492
rect 1582 488 1586 492
rect 1814 488 1818 492
rect 1910 488 1914 492
rect 142 478 146 482
rect 270 478 274 482
rect 390 478 394 482
rect 582 478 586 482
rect 678 478 682 482
rect 998 478 1002 482
rect 1030 478 1034 482
rect 1070 478 1074 482
rect 1190 478 1194 482
rect 1502 478 1506 482
rect 1510 478 1514 482
rect 1526 478 1530 482
rect 1686 478 1690 482
rect 1702 478 1706 482
rect 86 468 90 472
rect 158 468 162 472
rect 206 468 210 472
rect 382 468 386 472
rect 406 468 410 472
rect 454 468 458 472
rect 558 468 562 472
rect 638 468 642 472
rect 734 468 738 472
rect 806 468 810 472
rect 814 468 818 472
rect 878 468 882 472
rect 902 468 906 472
rect 926 468 930 472
rect 1078 468 1082 472
rect 1134 468 1138 472
rect 1278 468 1282 472
rect 1446 468 1450 472
rect 1526 468 1530 472
rect 1662 468 1666 472
rect 1694 468 1698 472
rect 1734 468 1738 472
rect 22 458 26 462
rect 94 459 98 463
rect 126 458 130 462
rect 142 458 146 462
rect 182 458 186 462
rect 278 458 282 462
rect 302 458 306 462
rect 422 458 426 462
rect 542 459 546 463
rect 742 458 746 462
rect 990 458 994 462
rect 1030 458 1034 462
rect 1086 458 1090 462
rect 1158 458 1162 462
rect 1262 459 1266 463
rect 1326 458 1330 462
rect 1454 459 1458 463
rect 1518 458 1522 462
rect 1542 458 1546 462
rect 1566 458 1570 462
rect 1646 459 1650 463
rect 1702 458 1706 462
rect 1718 458 1722 462
rect 1750 459 1754 463
rect 1854 458 1858 462
rect 1870 458 1874 462
rect 1918 458 1922 462
rect 782 448 786 452
rect 830 448 834 452
rect 846 448 850 452
rect 902 448 906 452
rect 918 448 922 452
rect 1574 448 1578 452
rect 1678 448 1682 452
rect 6 438 10 442
rect 1214 438 1218 442
rect 1558 438 1562 442
rect 1598 438 1602 442
rect 478 418 482 422
rect 458 403 462 407
rect 465 403 469 407
rect 1482 403 1486 407
rect 1489 403 1493 407
rect 6 388 10 392
rect 102 388 106 392
rect 286 388 290 392
rect 430 388 434 392
rect 534 388 538 392
rect 886 388 890 392
rect 982 388 986 392
rect 998 388 1002 392
rect 1246 388 1250 392
rect 1446 388 1450 392
rect 1566 388 1570 392
rect 1662 388 1666 392
rect 782 368 786 372
rect 1126 368 1130 372
rect 1350 368 1354 372
rect 1870 368 1874 372
rect 1902 368 1906 372
rect 70 347 74 351
rect 142 348 146 352
rect 222 347 226 351
rect 358 347 362 351
rect 398 348 402 352
rect 430 348 434 352
rect 446 348 450 352
rect 494 348 498 352
rect 510 348 514 352
rect 526 348 530 352
rect 574 348 578 352
rect 86 338 90 342
rect 238 338 242 342
rect 390 338 394 342
rect 598 347 602 351
rect 694 348 698 352
rect 1142 358 1146 362
rect 846 348 850 352
rect 918 347 922 351
rect 1062 348 1066 352
rect 1102 348 1106 352
rect 1190 347 1194 351
rect 1238 348 1242 352
rect 1302 348 1306 352
rect 1358 348 1362 352
rect 1510 348 1514 352
rect 1622 348 1626 352
rect 1678 348 1682 352
rect 1734 348 1738 352
rect 1758 348 1762 352
rect 1822 347 1826 351
rect 1894 348 1898 352
rect 1918 348 1922 352
rect 502 338 506 342
rect 542 338 546 342
rect 614 338 618 342
rect 678 338 682 342
rect 718 338 722 342
rect 750 338 754 342
rect 838 338 842 342
rect 1022 340 1026 344
rect 1030 338 1034 342
rect 1046 338 1050 342
rect 1206 338 1210 342
rect 1294 338 1298 342
rect 1390 338 1394 342
rect 1582 338 1586 342
rect 1686 338 1690 342
rect 326 328 330 332
rect 358 328 362 332
rect 526 328 530 332
rect 654 328 658 332
rect 662 328 666 332
rect 678 328 682 332
rect 758 328 762 332
rect 782 328 786 332
rect 918 328 922 332
rect 1046 328 1050 332
rect 1102 328 1106 332
rect 1118 328 1122 332
rect 1222 328 1226 332
rect 1502 328 1506 332
rect 1670 328 1674 332
rect 1926 327 1930 331
rect 294 318 298 322
rect 1054 318 1058 322
rect 1446 318 1450 322
rect 1702 318 1706 322
rect 1886 318 1890 322
rect 970 303 974 307
rect 977 303 981 307
rect 366 288 370 292
rect 382 288 386 292
rect 486 288 490 292
rect 542 288 546 292
rect 1222 288 1226 292
rect 1238 288 1242 292
rect 1542 288 1546 292
rect 1646 288 1650 292
rect 1678 288 1682 292
rect 1782 288 1786 292
rect 1886 288 1890 292
rect 6 278 10 282
rect 70 278 74 282
rect 142 278 146 282
rect 390 278 394 282
rect 686 278 690 282
rect 694 278 698 282
rect 718 278 722 282
rect 1054 278 1058 282
rect 1086 278 1090 282
rect 1182 278 1186 282
rect 1622 278 1626 282
rect 1774 278 1778 282
rect 1902 279 1906 283
rect 38 268 42 272
rect 94 268 98 272
rect 286 268 290 272
rect 406 268 410 272
rect 510 268 514 272
rect 598 268 602 272
rect 766 268 770 272
rect 838 268 842 272
rect 918 268 922 272
rect 958 268 962 272
rect 990 268 994 272
rect 1294 268 1298 272
rect 1350 268 1354 272
rect 1446 268 1450 272
rect 1670 268 1674 272
rect 1686 268 1690 272
rect 1806 268 1810 272
rect 118 258 122 262
rect 206 259 210 263
rect 238 258 242 262
rect 302 259 306 263
rect 374 258 378 262
rect 422 259 426 263
rect 606 259 610 263
rect 654 258 658 262
rect 718 258 722 262
rect 742 258 746 262
rect 766 258 770 262
rect 846 259 850 263
rect 934 258 938 262
rect 1086 259 1090 263
rect 1174 258 1178 262
rect 1334 258 1338 262
rect 1374 258 1378 262
rect 1486 258 1490 262
rect 1574 259 1578 263
rect 1598 258 1602 262
rect 1710 258 1714 262
rect 1742 259 1746 263
rect 1790 258 1794 262
rect 1822 259 1826 263
rect 1910 258 1914 262
rect 1918 258 1922 262
rect 734 248 738 252
rect 1646 248 1650 252
rect 70 238 74 242
rect 742 238 746 242
rect 750 238 754 242
rect 1134 238 1138 242
rect 1414 238 1418 242
rect 1926 238 1930 242
rect 174 218 178 222
rect 270 218 274 222
rect 782 218 786 222
rect 878 218 882 222
rect 1022 218 1026 222
rect 1118 218 1122 222
rect 1238 218 1242 222
rect 1430 218 1434 222
rect 1886 218 1890 222
rect 458 203 462 207
rect 465 203 469 207
rect 1482 203 1486 207
rect 1489 203 1493 207
rect 254 188 258 192
rect 598 188 602 192
rect 814 188 818 192
rect 878 188 882 192
rect 918 188 922 192
rect 1110 188 1114 192
rect 1526 188 1530 192
rect 1742 188 1746 192
rect 1846 188 1850 192
rect 350 168 354 172
rect 366 168 370 172
rect 494 168 498 172
rect 758 168 762 172
rect 1502 168 1506 172
rect 318 158 322 162
rect 782 158 786 162
rect 886 158 890 162
rect 1062 158 1066 162
rect 1094 158 1098 162
rect 1334 158 1338 162
rect 1390 158 1394 162
rect 1686 158 1690 162
rect 1758 158 1762 162
rect 1782 158 1786 162
rect 22 148 26 152
rect 86 148 90 152
rect 126 148 130 152
rect 174 147 178 151
rect 206 148 210 152
rect 246 148 250 152
rect 270 148 274 152
rect 342 148 346 152
rect 406 148 410 152
rect 470 148 474 152
rect 550 148 554 152
rect 694 148 698 152
rect 774 148 778 152
rect 814 148 818 152
rect 902 148 906 152
rect 918 148 922 152
rect 942 148 946 152
rect 1006 148 1010 152
rect 1150 148 1154 152
rect 1174 148 1178 152
rect 1190 148 1194 152
rect 1246 148 1250 152
rect 6 138 10 142
rect 110 138 114 142
rect 278 138 282 142
rect 302 138 306 142
rect 430 138 434 142
rect 462 138 466 142
rect 574 138 578 142
rect 590 138 594 142
rect 654 138 658 142
rect 670 138 674 142
rect 790 138 794 142
rect 806 138 810 142
rect 862 138 866 142
rect 910 138 914 142
rect 990 138 994 142
rect 1038 138 1042 142
rect 1070 138 1074 142
rect 1278 147 1282 151
rect 1350 148 1354 152
rect 1374 148 1378 152
rect 1390 148 1394 152
rect 1398 148 1402 152
rect 1358 138 1362 142
rect 1366 138 1370 142
rect 1454 147 1458 151
rect 1558 148 1562 152
rect 1630 148 1634 152
rect 1710 148 1714 152
rect 1734 148 1738 152
rect 1790 148 1794 152
rect 1798 148 1802 152
rect 1814 148 1818 152
rect 1830 148 1834 152
rect 1878 147 1882 151
rect 1406 138 1410 142
rect 1542 138 1546 142
rect 1574 138 1578 142
rect 1582 138 1586 142
rect 1702 138 1706 142
rect 1774 138 1778 142
rect 1806 138 1810 142
rect 1862 138 1866 142
rect 14 127 18 131
rect 142 128 146 132
rect 262 128 266 132
rect 286 128 290 132
rect 294 128 298 132
rect 310 128 314 132
rect 342 128 346 132
rect 798 128 802 132
rect 830 128 834 132
rect 838 128 842 132
rect 934 128 938 132
rect 950 127 954 131
rect 1006 128 1010 132
rect 1118 128 1122 132
rect 1230 128 1234 132
rect 1310 128 1314 132
rect 1422 128 1426 132
rect 1454 128 1458 132
rect 1550 128 1554 132
rect 1582 128 1586 132
rect 1830 128 1834 132
rect 1838 128 1842 132
rect 30 118 34 122
rect 134 118 138 122
rect 238 118 242 122
rect 486 118 490 122
rect 750 118 754 122
rect 998 118 1002 122
rect 1054 118 1058 122
rect 1158 118 1162 122
rect 1318 118 1322 122
rect 1414 118 1418 122
rect 1678 118 1682 122
rect 1686 118 1690 122
rect 1758 118 1762 122
rect 1942 118 1946 122
rect 970 103 974 107
rect 977 103 981 107
rect 118 88 122 92
rect 190 88 194 92
rect 302 88 306 92
rect 334 88 338 92
rect 350 88 354 92
rect 502 88 506 92
rect 638 88 642 92
rect 774 88 778 92
rect 814 88 818 92
rect 870 88 874 92
rect 1030 88 1034 92
rect 1054 88 1058 92
rect 1182 88 1186 92
rect 1374 88 1378 92
rect 1406 88 1410 92
rect 1502 88 1506 92
rect 1726 88 1730 92
rect 1942 88 1946 92
rect 6 78 10 82
rect 70 78 74 82
rect 126 78 130 82
rect 158 78 162 82
rect 174 78 178 82
rect 270 78 274 82
rect 302 78 306 82
rect 414 78 418 82
rect 494 78 498 82
rect 518 78 522 82
rect 574 79 578 83
rect 606 78 610 82
rect 614 78 618 82
rect 670 78 674 82
rect 742 78 746 82
rect 750 78 754 82
rect 782 78 786 82
rect 790 78 794 82
rect 822 78 826 82
rect 918 78 922 82
rect 1006 78 1010 82
rect 1214 78 1218 82
rect 1222 78 1226 82
rect 1438 78 1442 82
rect 1590 78 1594 82
rect 1622 78 1626 82
rect 1654 79 1658 83
rect 1822 78 1826 82
rect 1838 78 1842 82
rect 86 68 90 72
rect 118 68 122 72
rect 182 68 186 72
rect 214 68 218 72
rect 222 68 226 72
rect 238 68 242 72
rect 310 68 314 72
rect 462 68 466 72
rect 598 68 602 72
rect 622 68 626 72
rect 766 68 770 72
rect 798 68 802 72
rect 886 68 890 72
rect 1014 68 1018 72
rect 1046 68 1050 72
rect 1134 68 1138 72
rect 1198 68 1202 72
rect 1222 68 1226 72
rect 1246 68 1250 72
rect 1262 68 1266 72
rect 1294 68 1298 72
rect 1670 68 1674 72
rect 1718 68 1722 72
rect 1854 68 1858 72
rect 30 58 34 62
rect 142 58 146 62
rect 158 58 162 62
rect 206 58 210 62
rect 254 58 258 62
rect 294 58 298 62
rect 414 59 418 63
rect 454 58 458 62
rect 494 58 498 62
rect 510 58 514 62
rect 534 58 538 62
rect 566 58 570 62
rect 590 58 594 62
rect 694 58 698 62
rect 854 58 858 62
rect 926 58 930 62
rect 1022 58 1026 62
rect 1070 58 1074 62
rect 1150 59 1154 63
rect 1182 58 1186 62
rect 1206 58 1210 62
rect 1230 58 1234 62
rect 1262 58 1266 62
rect 1318 58 1322 62
rect 1390 58 1394 62
rect 1446 58 1450 62
rect 1582 58 1586 62
rect 1638 58 1642 62
rect 1646 58 1650 62
rect 1670 58 1674 62
rect 1718 58 1722 62
rect 1758 58 1762 62
rect 1782 58 1786 62
rect 1822 58 1826 62
rect 1878 58 1882 62
rect 46 48 50 52
rect 166 48 170 52
rect 190 48 194 52
rect 326 48 330 52
rect 486 48 490 52
rect 542 48 546 52
rect 558 48 562 52
rect 638 48 642 52
rect 870 48 874 52
rect 1030 48 1034 52
rect 1254 48 1258 52
rect 1278 48 1282 52
rect 1630 48 1634 52
rect 1694 48 1698 52
rect 854 38 858 42
rect 982 38 986 42
rect 1086 38 1090 42
rect 846 28 850 32
rect 582 18 586 22
rect 458 3 462 7
rect 465 3 469 7
rect 1482 3 1486 7
rect 1489 3 1493 7
<< metal2 >>
rect 166 1731 170 1732
rect 214 1731 218 1732
rect 830 1731 834 1732
rect 878 1731 882 1732
rect 166 1728 177 1731
rect 214 1728 225 1731
rect 174 1692 177 1728
rect 222 1692 225 1728
rect 822 1728 834 1731
rect 870 1728 882 1731
rect 1062 1728 1066 1732
rect 1078 1728 1082 1732
rect 1094 1731 1098 1732
rect 1094 1728 1105 1731
rect 822 1692 825 1728
rect 870 1692 873 1728
rect 968 1703 970 1707
rect 974 1703 977 1707
rect 981 1703 984 1707
rect 1062 1702 1065 1728
rect 1078 1692 1081 1728
rect 202 1678 206 1681
rect 426 1678 430 1681
rect 1046 1679 1054 1681
rect 1062 1682 1065 1688
rect 1046 1678 1057 1679
rect 6 1672 9 1678
rect 62 1672 65 1678
rect 22 1662 25 1668
rect 30 1652 33 1668
rect 54 1662 57 1668
rect 70 1642 73 1678
rect 94 1672 97 1678
rect 114 1668 118 1671
rect 82 1658 86 1661
rect 102 1642 105 1658
rect 118 1652 121 1658
rect 126 1592 129 1678
rect 134 1672 137 1678
rect 142 1642 145 1668
rect 182 1662 185 1668
rect 162 1658 166 1661
rect 150 1652 153 1658
rect 6 1442 9 1518
rect 62 1472 65 1548
rect 62 1462 65 1468
rect 10 1438 14 1441
rect 70 1402 73 1528
rect 6 1362 9 1368
rect 62 1342 65 1348
rect 70 1342 73 1398
rect 62 1262 65 1298
rect 10 1238 14 1241
rect 6 1192 9 1238
rect 62 1152 65 1258
rect 70 1142 73 1338
rect 86 1282 89 1468
rect 102 1451 105 1548
rect 142 1542 145 1548
rect 150 1542 153 1648
rect 214 1592 217 1678
rect 406 1672 409 1678
rect 294 1652 297 1659
rect 234 1618 238 1621
rect 254 1552 257 1618
rect 262 1592 265 1638
rect 310 1572 313 1668
rect 390 1652 393 1659
rect 322 1618 326 1621
rect 202 1548 206 1551
rect 358 1551 361 1558
rect 110 1462 113 1468
rect 118 1462 121 1468
rect 146 1458 150 1461
rect 102 1448 113 1451
rect 86 1272 89 1278
rect 110 1272 113 1448
rect 126 1352 129 1458
rect 134 1442 137 1458
rect 158 1372 161 1548
rect 166 1462 169 1548
rect 190 1542 193 1548
rect 206 1512 209 1548
rect 238 1542 241 1548
rect 238 1463 241 1478
rect 254 1462 257 1548
rect 286 1542 289 1548
rect 374 1542 377 1558
rect 298 1518 302 1521
rect 178 1418 182 1421
rect 134 1342 137 1348
rect 142 1332 145 1338
rect 142 1272 145 1328
rect 158 1262 161 1368
rect 190 1362 193 1368
rect 198 1342 201 1348
rect 206 1332 209 1458
rect 254 1421 257 1458
rect 254 1418 265 1421
rect 230 1352 233 1358
rect 214 1332 217 1348
rect 222 1342 225 1348
rect 194 1328 198 1331
rect 166 1263 169 1268
rect 86 1082 89 1238
rect 102 1172 105 1218
rect 122 1148 126 1151
rect 134 1144 137 1148
rect 122 1138 126 1141
rect 138 1140 142 1143
rect 134 1138 137 1140
rect 102 1132 105 1138
rect 182 1132 185 1268
rect 190 1132 193 1148
rect 110 1092 113 1118
rect 150 1082 153 1118
rect 74 1078 78 1081
rect 10 1068 14 1071
rect 86 1070 89 1078
rect 110 1072 113 1078
rect 22 1042 25 1048
rect 54 1042 57 1058
rect 26 958 30 961
rect 6 942 9 948
rect 14 892 17 958
rect 54 952 57 1038
rect 26 948 30 951
rect 10 868 14 871
rect 22 852 25 898
rect 38 862 41 908
rect 54 902 57 948
rect 78 942 81 1068
rect 126 1062 129 1078
rect 134 1062 137 1068
rect 158 1062 161 1088
rect 166 1072 169 1078
rect 174 1072 177 1078
rect 106 1058 110 1061
rect 142 1052 145 1058
rect 126 1042 129 1048
rect 154 1018 158 1021
rect 138 988 142 991
rect 62 938 70 941
rect 62 872 65 938
rect 126 932 129 938
rect 74 928 78 931
rect 106 918 110 921
rect 62 862 65 868
rect 86 862 89 918
rect 118 862 121 908
rect 126 892 129 928
rect 54 752 57 818
rect 62 792 65 858
rect 78 852 81 858
rect 102 802 105 818
rect 98 788 102 791
rect 74 748 78 751
rect 6 742 9 748
rect 94 742 97 748
rect 74 738 78 741
rect 22 662 25 708
rect 30 672 33 738
rect 94 672 97 728
rect 102 692 105 718
rect 6 642 9 648
rect 30 632 33 668
rect 30 542 33 628
rect 10 538 14 541
rect 86 531 89 618
rect 94 552 97 568
rect 102 552 105 558
rect 110 542 113 548
rect 82 528 89 531
rect 22 462 25 508
rect 34 488 38 491
rect 6 442 9 448
rect 10 388 14 391
rect 62 302 65 518
rect 86 482 89 528
rect 86 472 89 478
rect 70 351 73 358
rect 86 342 89 468
rect 94 463 97 528
rect 110 492 113 538
rect 118 491 121 798
rect 126 562 129 568
rect 134 552 137 898
rect 166 822 169 948
rect 182 942 185 1128
rect 230 1071 233 1348
rect 242 1328 246 1331
rect 238 1262 241 1318
rect 254 1262 257 1398
rect 262 1352 265 1418
rect 270 1362 273 1418
rect 286 1402 289 1438
rect 298 1348 302 1351
rect 270 1331 273 1348
rect 310 1332 313 1498
rect 326 1472 329 1538
rect 414 1511 417 1547
rect 406 1508 417 1511
rect 422 1542 425 1678
rect 622 1672 625 1678
rect 430 1662 433 1668
rect 438 1662 441 1668
rect 574 1663 577 1668
rect 482 1658 486 1661
rect 618 1658 622 1661
rect 666 1658 670 1661
rect 446 1582 449 1658
rect 470 1622 473 1658
rect 494 1652 497 1658
rect 514 1618 518 1621
rect 456 1603 458 1607
rect 462 1603 465 1607
rect 469 1603 472 1607
rect 550 1562 553 1658
rect 606 1642 609 1658
rect 550 1552 553 1558
rect 406 1492 409 1508
rect 422 1502 425 1538
rect 510 1532 513 1538
rect 474 1518 478 1521
rect 334 1463 337 1478
rect 398 1472 401 1478
rect 430 1472 433 1518
rect 510 1502 513 1528
rect 522 1518 526 1521
rect 566 1512 569 1588
rect 574 1512 577 1548
rect 598 1532 601 1538
rect 610 1518 614 1521
rect 534 1482 537 1488
rect 370 1468 374 1471
rect 426 1468 430 1471
rect 514 1468 518 1471
rect 378 1458 382 1461
rect 370 1448 374 1451
rect 358 1352 361 1388
rect 366 1362 369 1448
rect 390 1442 393 1468
rect 414 1462 417 1468
rect 422 1442 425 1458
rect 382 1372 385 1428
rect 342 1348 350 1351
rect 318 1342 321 1348
rect 326 1342 329 1348
rect 270 1328 278 1331
rect 302 1322 305 1328
rect 342 1312 345 1348
rect 286 1292 289 1308
rect 302 1282 305 1288
rect 334 1272 337 1278
rect 306 1268 310 1271
rect 294 1262 297 1268
rect 330 1258 334 1261
rect 254 1152 257 1258
rect 342 1251 345 1278
rect 338 1248 345 1251
rect 334 1242 337 1248
rect 286 1172 289 1218
rect 286 1152 289 1158
rect 350 1152 353 1338
rect 366 1231 369 1358
rect 382 1352 385 1368
rect 390 1342 393 1438
rect 422 1352 425 1438
rect 438 1431 441 1468
rect 526 1462 529 1468
rect 566 1462 569 1508
rect 582 1472 585 1518
rect 630 1511 633 1618
rect 630 1508 641 1511
rect 614 1492 617 1508
rect 626 1478 630 1481
rect 610 1468 617 1471
rect 574 1462 577 1468
rect 450 1458 454 1461
rect 430 1428 441 1431
rect 430 1362 433 1428
rect 438 1362 441 1418
rect 456 1403 458 1407
rect 462 1403 465 1407
rect 469 1403 472 1407
rect 510 1392 513 1458
rect 518 1442 521 1458
rect 554 1448 558 1451
rect 518 1402 521 1438
rect 574 1402 577 1458
rect 542 1392 545 1398
rect 450 1368 457 1371
rect 418 1338 422 1341
rect 374 1332 377 1338
rect 394 1328 398 1331
rect 374 1272 377 1308
rect 406 1302 409 1318
rect 430 1312 433 1358
rect 438 1332 441 1338
rect 382 1272 385 1278
rect 374 1252 377 1258
rect 366 1228 377 1231
rect 354 1148 358 1151
rect 318 1132 321 1147
rect 354 1138 358 1141
rect 254 1112 257 1118
rect 238 1082 241 1088
rect 294 1072 297 1078
rect 230 1068 238 1071
rect 302 1062 305 1068
rect 346 1058 350 1061
rect 222 1052 225 1058
rect 318 1052 321 1058
rect 194 1048 198 1051
rect 190 1042 193 1048
rect 222 1001 225 1048
rect 222 998 233 1001
rect 194 947 198 950
rect 150 742 153 818
rect 162 748 166 751
rect 146 738 150 741
rect 166 663 169 748
rect 182 672 185 868
rect 190 863 193 947
rect 230 892 233 998
rect 262 952 265 1018
rect 270 942 273 1018
rect 318 982 321 1048
rect 282 948 286 951
rect 310 942 313 948
rect 258 938 262 941
rect 298 928 302 931
rect 270 922 273 928
rect 318 912 321 978
rect 358 972 361 1138
rect 366 1092 369 1218
rect 374 1162 377 1228
rect 374 1091 377 1158
rect 382 1102 385 1268
rect 422 1262 425 1278
rect 398 1252 401 1258
rect 430 1252 433 1288
rect 438 1272 441 1278
rect 446 1261 449 1348
rect 454 1292 457 1368
rect 558 1342 561 1348
rect 566 1342 569 1358
rect 478 1292 481 1338
rect 438 1258 449 1261
rect 486 1262 489 1288
rect 494 1272 497 1335
rect 526 1322 529 1338
rect 510 1292 513 1298
rect 518 1282 521 1288
rect 526 1272 529 1278
rect 526 1262 529 1268
rect 394 1238 398 1241
rect 410 1238 414 1241
rect 422 1232 425 1248
rect 438 1192 441 1258
rect 502 1252 505 1258
rect 456 1203 458 1207
rect 462 1203 465 1207
rect 469 1203 472 1207
rect 398 1142 401 1178
rect 426 1168 430 1171
rect 442 1168 446 1171
rect 478 1162 481 1198
rect 490 1168 494 1171
rect 502 1162 505 1218
rect 518 1182 521 1188
rect 514 1168 518 1171
rect 522 1168 526 1171
rect 542 1162 545 1318
rect 554 1258 558 1261
rect 558 1242 561 1248
rect 550 1212 553 1218
rect 566 1202 569 1308
rect 574 1302 577 1348
rect 582 1291 585 1468
rect 594 1458 598 1461
rect 590 1362 593 1418
rect 614 1392 617 1468
rect 638 1462 641 1508
rect 646 1492 649 1638
rect 670 1512 673 1548
rect 694 1542 697 1668
rect 726 1622 729 1648
rect 726 1562 729 1618
rect 694 1532 697 1538
rect 710 1512 713 1518
rect 686 1492 689 1498
rect 710 1482 713 1488
rect 630 1442 633 1458
rect 630 1392 633 1438
rect 638 1432 641 1458
rect 662 1412 665 1458
rect 670 1392 673 1468
rect 726 1462 729 1558
rect 774 1542 777 1547
rect 774 1472 777 1528
rect 702 1382 705 1458
rect 714 1448 718 1451
rect 734 1432 737 1468
rect 746 1418 750 1421
rect 782 1392 785 1468
rect 790 1461 793 1659
rect 806 1632 809 1668
rect 822 1572 825 1628
rect 846 1542 849 1678
rect 866 1658 870 1661
rect 890 1658 894 1661
rect 806 1512 809 1518
rect 870 1511 873 1547
rect 870 1508 881 1511
rect 878 1492 881 1508
rect 842 1478 846 1481
rect 822 1472 825 1478
rect 886 1472 889 1538
rect 902 1532 905 1678
rect 974 1663 977 1668
rect 1010 1658 1014 1661
rect 942 1632 945 1658
rect 1022 1652 1025 1678
rect 1046 1662 1049 1678
rect 1038 1652 1041 1658
rect 914 1618 918 1621
rect 1074 1618 1078 1621
rect 1102 1621 1105 1728
rect 1158 1728 1162 1732
rect 1174 1731 1178 1732
rect 1166 1728 1178 1731
rect 1198 1731 1202 1732
rect 1198 1728 1209 1731
rect 1158 1702 1161 1728
rect 1166 1692 1169 1728
rect 1206 1692 1209 1728
rect 1310 1728 1314 1732
rect 1326 1728 1330 1732
rect 1342 1731 1346 1732
rect 1342 1728 1353 1731
rect 1310 1692 1313 1728
rect 1326 1702 1329 1728
rect 1350 1692 1353 1728
rect 1510 1728 1514 1732
rect 1678 1728 1682 1732
rect 1702 1728 1706 1732
rect 1742 1731 1746 1732
rect 1758 1731 1762 1732
rect 1862 1731 1866 1732
rect 1742 1728 1753 1731
rect 1758 1728 1769 1731
rect 1510 1702 1513 1728
rect 1450 1678 1454 1681
rect 1150 1672 1153 1678
rect 1382 1672 1385 1678
rect 1510 1672 1513 1678
rect 1270 1662 1273 1668
rect 1122 1658 1126 1661
rect 1094 1618 1105 1621
rect 1070 1592 1073 1608
rect 1094 1592 1097 1618
rect 986 1568 990 1571
rect 1018 1558 1022 1561
rect 910 1552 913 1558
rect 950 1552 953 1558
rect 1030 1552 1033 1568
rect 1110 1552 1113 1618
rect 1118 1592 1121 1648
rect 1150 1592 1153 1658
rect 1182 1562 1185 1658
rect 1190 1602 1193 1658
rect 1246 1632 1249 1658
rect 1326 1641 1329 1658
rect 1322 1638 1329 1641
rect 1214 1582 1217 1618
rect 1270 1592 1273 1598
rect 1238 1552 1241 1558
rect 1286 1552 1289 1558
rect 1294 1552 1297 1598
rect 1318 1592 1321 1628
rect 1002 1548 1006 1551
rect 1018 1548 1022 1551
rect 1082 1548 1086 1551
rect 1218 1548 1222 1551
rect 1258 1548 1262 1551
rect 926 1532 929 1538
rect 866 1468 870 1471
rect 790 1459 798 1461
rect 802 1459 806 1462
rect 838 1462 841 1468
rect 910 1462 913 1488
rect 918 1462 921 1468
rect 942 1462 945 1548
rect 950 1492 953 1548
rect 958 1542 961 1548
rect 970 1528 974 1531
rect 1042 1528 1046 1531
rect 968 1503 970 1507
rect 974 1503 977 1507
rect 981 1503 984 1507
rect 1014 1492 1017 1528
rect 1042 1488 1046 1491
rect 790 1458 801 1459
rect 866 1458 870 1461
rect 854 1442 857 1458
rect 638 1362 641 1378
rect 650 1368 662 1371
rect 682 1368 689 1371
rect 662 1362 665 1368
rect 590 1342 593 1358
rect 614 1352 617 1358
rect 630 1352 633 1358
rect 618 1338 622 1341
rect 574 1288 585 1291
rect 574 1282 577 1288
rect 594 1278 598 1281
rect 566 1162 569 1198
rect 554 1158 558 1161
rect 454 1152 457 1158
rect 498 1148 502 1151
rect 406 1142 409 1148
rect 390 1122 393 1128
rect 374 1088 385 1091
rect 370 1078 374 1081
rect 370 1068 374 1071
rect 350 962 353 968
rect 334 952 337 958
rect 358 942 361 968
rect 374 952 377 1038
rect 382 962 385 1088
rect 398 1052 401 1098
rect 406 1062 409 1078
rect 414 1072 417 1128
rect 430 1082 433 1148
rect 510 1142 513 1158
rect 538 1148 542 1151
rect 574 1141 577 1278
rect 614 1272 617 1338
rect 638 1312 641 1348
rect 654 1322 657 1338
rect 654 1292 657 1318
rect 662 1281 665 1358
rect 674 1348 678 1351
rect 686 1322 689 1368
rect 738 1368 742 1371
rect 710 1362 713 1368
rect 718 1362 721 1368
rect 710 1352 713 1358
rect 806 1352 809 1438
rect 814 1352 817 1418
rect 830 1392 833 1438
rect 862 1432 865 1458
rect 890 1448 894 1451
rect 886 1362 889 1448
rect 902 1412 905 1428
rect 694 1342 697 1348
rect 726 1342 729 1348
rect 738 1338 742 1341
rect 654 1278 665 1281
rect 614 1252 617 1268
rect 630 1252 633 1258
rect 586 1238 590 1241
rect 598 1162 601 1248
rect 594 1158 598 1161
rect 626 1158 630 1161
rect 586 1148 590 1151
rect 574 1138 582 1141
rect 510 1112 513 1138
rect 570 1128 574 1131
rect 390 1042 393 1048
rect 398 992 401 1048
rect 406 1032 409 1048
rect 418 1038 422 1041
rect 394 948 398 951
rect 330 938 334 941
rect 342 932 345 938
rect 270 892 273 908
rect 342 892 345 918
rect 366 902 369 948
rect 382 942 385 948
rect 414 942 417 958
rect 430 951 433 1068
rect 446 972 449 1078
rect 462 1042 465 1088
rect 550 1062 553 1068
rect 574 1062 577 1118
rect 474 1058 478 1061
rect 534 1022 537 1058
rect 456 1003 458 1007
rect 462 1003 465 1007
rect 469 1003 472 1007
rect 518 952 521 1018
rect 542 1012 545 1058
rect 422 948 433 951
rect 466 948 470 951
rect 390 932 393 938
rect 398 892 401 938
rect 422 922 425 948
rect 478 942 481 948
rect 534 942 537 968
rect 542 962 545 978
rect 558 962 561 1018
rect 434 938 438 941
rect 462 932 465 938
rect 434 928 438 931
rect 322 878 326 881
rect 282 868 286 871
rect 230 722 233 748
rect 238 682 241 868
rect 302 862 305 868
rect 254 832 257 858
rect 182 662 185 668
rect 158 592 161 648
rect 198 642 201 648
rect 222 622 225 658
rect 182 592 185 618
rect 254 572 257 828
rect 286 792 289 818
rect 318 792 321 878
rect 350 872 353 878
rect 382 872 385 878
rect 362 868 366 871
rect 354 848 358 851
rect 318 772 321 788
rect 310 752 313 758
rect 290 728 294 731
rect 166 542 169 558
rect 198 552 201 568
rect 230 552 233 558
rect 222 542 225 548
rect 146 538 150 541
rect 238 532 241 548
rect 246 532 249 538
rect 118 488 129 491
rect 126 462 129 488
rect 138 478 142 481
rect 158 472 161 478
rect 182 462 185 498
rect 206 472 209 528
rect 214 502 217 518
rect 238 492 241 528
rect 270 482 273 668
rect 302 661 305 718
rect 298 658 305 661
rect 278 552 281 638
rect 286 592 289 648
rect 294 562 297 618
rect 318 562 321 718
rect 334 692 337 818
rect 342 812 345 848
rect 366 742 369 868
rect 378 848 382 851
rect 390 792 393 868
rect 406 852 409 898
rect 446 892 449 918
rect 454 882 457 888
rect 442 878 446 881
rect 442 868 446 871
rect 470 862 473 938
rect 558 922 561 938
rect 486 872 489 918
rect 518 892 521 898
rect 534 872 537 878
rect 426 858 430 861
rect 462 852 465 858
rect 414 842 417 848
rect 430 842 433 848
rect 422 792 425 808
rect 456 803 458 807
rect 462 803 465 807
rect 469 803 472 807
rect 454 762 457 768
rect 430 752 433 758
rect 478 752 481 868
rect 542 852 545 918
rect 566 862 569 978
rect 582 952 585 1138
rect 606 1132 609 1148
rect 614 1142 617 1148
rect 630 1132 633 1138
rect 638 1131 641 1268
rect 654 1242 657 1278
rect 662 1268 678 1271
rect 662 1262 665 1268
rect 694 1262 697 1338
rect 710 1332 713 1338
rect 750 1332 753 1338
rect 670 1252 673 1258
rect 678 1252 681 1258
rect 670 1232 673 1248
rect 694 1192 697 1228
rect 654 1152 657 1168
rect 686 1152 689 1168
rect 710 1152 713 1328
rect 718 1292 721 1318
rect 726 1282 729 1288
rect 718 1272 721 1278
rect 726 1252 729 1258
rect 766 1232 769 1278
rect 782 1272 785 1335
rect 798 1272 801 1338
rect 798 1262 801 1268
rect 798 1242 801 1248
rect 778 1238 782 1241
rect 758 1151 761 1178
rect 774 1132 777 1138
rect 798 1132 801 1168
rect 806 1162 809 1348
rect 814 1202 817 1348
rect 838 1322 841 1348
rect 846 1342 849 1348
rect 854 1342 857 1348
rect 838 1302 841 1318
rect 826 1288 830 1291
rect 838 1272 841 1278
rect 826 1248 830 1251
rect 838 1172 841 1268
rect 870 1262 873 1318
rect 886 1312 889 1358
rect 902 1352 905 1408
rect 878 1292 881 1308
rect 850 1258 854 1261
rect 870 1182 873 1258
rect 886 1252 889 1258
rect 838 1152 841 1158
rect 862 1152 865 1158
rect 814 1142 817 1148
rect 634 1128 641 1131
rect 614 1072 617 1078
rect 590 1062 593 1068
rect 622 1062 625 1108
rect 594 1048 598 1051
rect 606 1042 609 1048
rect 606 982 609 1038
rect 622 952 625 1018
rect 594 948 598 951
rect 574 902 577 938
rect 614 932 617 948
rect 630 942 633 1128
rect 670 1122 673 1128
rect 638 1082 641 1118
rect 662 1092 665 1118
rect 678 1112 681 1118
rect 646 1072 649 1078
rect 654 1072 657 1078
rect 674 1068 678 1071
rect 686 1070 689 1128
rect 766 1092 769 1098
rect 826 1088 830 1091
rect 838 1091 841 1148
rect 858 1138 862 1141
rect 854 1122 857 1138
rect 870 1102 873 1148
rect 894 1112 897 1148
rect 902 1102 905 1348
rect 918 1342 921 1458
rect 934 1432 937 1458
rect 942 1392 945 1448
rect 966 1352 969 1458
rect 930 1348 934 1351
rect 914 1338 918 1341
rect 968 1303 970 1307
rect 974 1303 977 1307
rect 981 1303 984 1307
rect 990 1272 993 1458
rect 1006 1352 1009 1378
rect 1014 1352 1017 1358
rect 962 1258 966 1261
rect 910 1232 913 1238
rect 982 1132 985 1138
rect 930 1128 934 1131
rect 870 1092 873 1098
rect 838 1088 849 1091
rect 702 1082 705 1088
rect 686 1062 689 1066
rect 750 1062 753 1078
rect 642 1058 646 1061
rect 658 1058 662 1061
rect 674 1058 678 1061
rect 706 1048 710 1051
rect 734 1042 737 1058
rect 774 1032 777 1078
rect 734 962 737 1008
rect 678 942 681 948
rect 630 932 633 938
rect 586 928 590 931
rect 582 912 585 918
rect 678 892 681 938
rect 686 932 689 938
rect 710 931 713 948
rect 710 928 721 931
rect 626 888 630 891
rect 582 882 585 888
rect 686 863 689 868
rect 602 858 606 861
rect 590 842 593 848
rect 598 792 601 838
rect 378 747 382 750
rect 374 672 377 738
rect 382 682 385 698
rect 338 648 342 651
rect 366 622 369 658
rect 370 618 377 621
rect 350 542 353 598
rect 374 562 377 618
rect 382 602 385 678
rect 398 672 401 728
rect 414 662 417 728
rect 422 712 425 748
rect 434 738 438 741
rect 474 728 478 731
rect 422 662 425 708
rect 486 692 489 768
rect 510 762 513 768
rect 558 762 561 768
rect 538 758 542 761
rect 518 751 521 758
rect 498 748 521 751
rect 602 748 606 751
rect 558 742 561 748
rect 566 742 569 748
rect 578 738 582 741
rect 534 732 537 738
rect 598 732 601 748
rect 614 742 617 818
rect 654 772 657 778
rect 638 768 646 771
rect 630 732 633 738
rect 498 728 502 731
rect 514 728 518 731
rect 526 682 529 718
rect 534 702 537 728
rect 502 662 505 678
rect 534 672 537 698
rect 550 672 553 678
rect 542 662 545 668
rect 566 662 569 668
rect 402 558 406 561
rect 278 532 281 538
rect 302 532 305 538
rect 358 532 361 558
rect 374 552 377 558
rect 422 532 425 538
rect 430 532 433 658
rect 534 652 537 658
rect 574 652 577 728
rect 598 672 601 718
rect 622 712 625 718
rect 630 692 633 698
rect 622 682 625 688
rect 638 682 641 768
rect 662 762 665 858
rect 654 752 657 758
rect 702 752 705 868
rect 718 852 721 928
rect 726 892 729 958
rect 734 952 737 958
rect 774 952 777 1028
rect 822 1002 825 1068
rect 806 952 809 958
rect 814 952 817 978
rect 838 952 841 1058
rect 846 952 849 1088
rect 894 1063 897 1088
rect 910 1072 913 1128
rect 918 1092 921 1118
rect 950 1112 953 1118
rect 942 1092 945 1098
rect 950 1092 953 1108
rect 968 1103 970 1107
rect 974 1103 977 1107
rect 981 1103 984 1107
rect 990 1072 993 1268
rect 1006 1252 1009 1348
rect 1030 1292 1033 1478
rect 1038 1392 1041 1478
rect 1070 1452 1073 1458
rect 1086 1392 1089 1528
rect 1102 1512 1105 1548
rect 1134 1492 1137 1548
rect 1102 1463 1105 1468
rect 1134 1362 1137 1418
rect 1150 1392 1153 1548
rect 1218 1538 1222 1541
rect 1194 1528 1198 1531
rect 1174 1482 1177 1528
rect 1198 1522 1201 1528
rect 1254 1522 1257 1538
rect 1278 1532 1281 1548
rect 1302 1542 1305 1548
rect 1234 1478 1238 1481
rect 1250 1478 1257 1481
rect 1214 1472 1217 1478
rect 1246 1472 1249 1478
rect 1254 1472 1257 1478
rect 1194 1459 1198 1462
rect 1234 1458 1241 1461
rect 1198 1392 1201 1428
rect 1238 1392 1241 1458
rect 1254 1352 1257 1358
rect 1262 1352 1265 1478
rect 1270 1352 1273 1508
rect 1278 1432 1281 1528
rect 1278 1352 1281 1418
rect 1294 1392 1297 1528
rect 1310 1382 1313 1578
rect 1382 1552 1385 1668
rect 1390 1662 1393 1668
rect 1454 1662 1457 1668
rect 1470 1662 1473 1668
rect 1526 1662 1529 1698
rect 1598 1662 1601 1668
rect 1506 1658 1510 1661
rect 1446 1622 1449 1658
rect 1494 1651 1497 1658
rect 1526 1652 1529 1658
rect 1494 1648 1505 1651
rect 1446 1582 1449 1618
rect 1480 1603 1482 1607
rect 1486 1603 1489 1607
rect 1493 1603 1496 1607
rect 1462 1552 1465 1558
rect 1478 1552 1481 1588
rect 1502 1552 1505 1648
rect 1546 1618 1550 1621
rect 1606 1572 1609 1668
rect 1618 1588 1622 1591
rect 1630 1581 1633 1638
rect 1622 1578 1633 1581
rect 1510 1552 1513 1558
rect 1402 1548 1406 1551
rect 1326 1532 1329 1548
rect 1342 1542 1345 1548
rect 1382 1532 1385 1548
rect 1326 1492 1329 1518
rect 1342 1472 1345 1528
rect 1350 1512 1353 1518
rect 1318 1442 1321 1468
rect 1390 1463 1393 1548
rect 1446 1542 1449 1548
rect 1454 1492 1457 1548
rect 1474 1488 1478 1491
rect 1486 1482 1489 1548
rect 1542 1542 1545 1548
rect 1526 1532 1529 1538
rect 1566 1532 1569 1548
rect 1514 1528 1518 1531
rect 1358 1452 1361 1458
rect 1422 1442 1425 1468
rect 1486 1462 1489 1478
rect 1518 1452 1521 1468
rect 1542 1462 1545 1528
rect 1606 1491 1609 1528
rect 1602 1488 1609 1491
rect 1622 1492 1625 1578
rect 1646 1552 1649 1648
rect 1670 1592 1673 1658
rect 1662 1552 1665 1558
rect 1662 1532 1665 1538
rect 1630 1482 1633 1518
rect 1670 1472 1673 1478
rect 1610 1468 1614 1471
rect 1678 1462 1681 1728
rect 1702 1702 1705 1728
rect 1686 1551 1689 1698
rect 1750 1692 1753 1728
rect 1694 1652 1697 1658
rect 1734 1641 1737 1658
rect 1734 1638 1742 1641
rect 1686 1548 1694 1551
rect 1694 1482 1697 1548
rect 1718 1532 1721 1548
rect 1726 1531 1729 1618
rect 1758 1582 1761 1618
rect 1758 1552 1761 1578
rect 1766 1562 1769 1728
rect 1854 1728 1866 1731
rect 1886 1731 1890 1732
rect 1910 1731 1914 1732
rect 1886 1728 1897 1731
rect 1910 1728 1921 1731
rect 1854 1692 1857 1728
rect 1894 1692 1897 1728
rect 1918 1692 1921 1728
rect 1866 1679 1873 1681
rect 1862 1678 1873 1679
rect 1794 1658 1798 1661
rect 1814 1592 1817 1658
rect 1794 1568 1801 1571
rect 1766 1552 1769 1558
rect 1798 1552 1801 1568
rect 1814 1552 1817 1588
rect 1722 1528 1729 1531
rect 1718 1482 1721 1488
rect 1734 1462 1737 1548
rect 1742 1542 1745 1548
rect 1774 1542 1777 1548
rect 1806 1542 1809 1548
rect 1822 1492 1825 1528
rect 1838 1521 1841 1668
rect 1870 1662 1873 1678
rect 1878 1641 1881 1658
rect 1878 1638 1886 1641
rect 1902 1641 1905 1658
rect 1926 1642 1929 1678
rect 1902 1638 1910 1641
rect 1914 1578 1918 1581
rect 1854 1551 1857 1558
rect 1926 1552 1929 1608
rect 1918 1548 1926 1551
rect 1830 1518 1841 1521
rect 1750 1482 1753 1488
rect 1830 1472 1833 1518
rect 1626 1458 1630 1461
rect 1626 1448 1630 1451
rect 1638 1432 1641 1458
rect 1702 1452 1705 1458
rect 1750 1452 1753 1459
rect 1658 1448 1662 1451
rect 1710 1442 1713 1448
rect 1322 1418 1326 1421
rect 1480 1403 1482 1407
rect 1486 1403 1489 1407
rect 1493 1403 1496 1407
rect 1614 1392 1617 1418
rect 1310 1352 1313 1378
rect 1498 1368 1502 1371
rect 1318 1362 1321 1368
rect 1374 1362 1377 1368
rect 1454 1362 1457 1368
rect 1546 1358 1550 1361
rect 1050 1348 1054 1351
rect 1234 1348 1238 1351
rect 1014 1122 1017 1147
rect 1030 1092 1033 1168
rect 1070 1152 1073 1348
rect 1102 1312 1105 1338
rect 1110 1332 1113 1348
rect 1102 1292 1105 1308
rect 1110 1292 1113 1328
rect 1090 1268 1094 1271
rect 1134 1262 1137 1348
rect 1174 1292 1177 1348
rect 1206 1322 1209 1348
rect 1174 1282 1177 1288
rect 1198 1282 1201 1288
rect 1226 1268 1230 1271
rect 1262 1262 1265 1348
rect 1270 1342 1273 1348
rect 1118 1242 1121 1258
rect 1102 1152 1105 1178
rect 1078 1142 1081 1148
rect 1034 1088 1038 1091
rect 1022 1072 1025 1078
rect 874 978 878 981
rect 910 952 913 1068
rect 994 1058 998 1061
rect 1070 1042 1073 1058
rect 718 822 721 848
rect 734 761 737 948
rect 742 892 745 948
rect 726 758 737 761
rect 774 762 777 948
rect 802 928 806 931
rect 814 922 817 948
rect 790 862 793 918
rect 846 892 849 948
rect 870 942 873 948
rect 910 932 913 948
rect 934 942 937 948
rect 990 942 993 998
rect 1030 992 1033 1018
rect 1046 992 1049 1038
rect 874 928 878 931
rect 878 891 881 918
rect 874 888 881 891
rect 702 722 705 748
rect 602 658 606 661
rect 590 652 593 658
rect 456 603 458 607
rect 462 603 465 607
rect 469 603 472 607
rect 446 552 449 558
rect 278 462 281 498
rect 302 492 305 528
rect 94 402 97 459
rect 98 388 102 391
rect 142 352 145 458
rect 222 351 225 398
rect 286 392 289 488
rect 302 462 305 478
rect 326 472 329 518
rect 430 502 433 528
rect 334 492 337 498
rect 382 492 385 498
rect 390 482 393 488
rect 406 472 409 498
rect 426 488 430 491
rect 454 472 457 558
rect 486 552 489 618
rect 510 562 513 578
rect 606 571 609 618
rect 598 568 609 571
rect 518 562 521 568
rect 494 542 497 558
rect 478 492 481 528
rect 482 488 486 491
rect 378 468 382 471
rect 286 362 289 388
rect 358 351 361 428
rect 406 392 409 468
rect 426 458 433 461
rect 430 392 433 458
rect 456 403 458 407
rect 462 403 465 407
rect 469 403 472 407
rect 478 362 481 418
rect 358 342 361 347
rect 390 342 393 358
rect 402 348 406 351
rect 450 348 454 351
rect 242 338 246 341
rect 86 291 89 338
rect 86 288 97 291
rect 6 252 9 278
rect 38 252 41 268
rect 70 252 73 278
rect 94 272 97 288
rect 74 238 78 241
rect 110 162 113 298
rect 142 272 145 278
rect 122 258 126 261
rect 238 262 241 338
rect 326 332 329 338
rect 298 318 302 321
rect 286 272 289 278
rect 206 252 209 259
rect 178 218 182 221
rect 6 142 9 148
rect 22 131 25 148
rect 18 128 25 131
rect 34 118 38 121
rect 6 82 9 118
rect 70 82 73 108
rect 86 72 89 148
rect 110 142 113 158
rect 126 102 129 148
rect 174 142 177 147
rect 142 122 145 128
rect 134 112 137 118
rect 122 88 126 91
rect 130 78 134 81
rect 170 78 174 81
rect 158 72 161 78
rect 182 72 185 218
rect 238 172 241 258
rect 302 232 305 259
rect 254 192 257 228
rect 266 218 270 221
rect 350 172 353 288
rect 358 271 361 328
rect 382 292 385 308
rect 366 282 369 288
rect 390 282 393 338
rect 406 272 409 278
rect 358 268 369 271
rect 366 172 369 268
rect 422 263 425 338
rect 430 312 433 348
rect 494 342 497 348
rect 502 342 505 358
rect 510 352 513 548
rect 578 547 582 550
rect 574 532 577 538
rect 558 472 561 478
rect 538 459 542 462
rect 530 388 534 391
rect 574 352 577 528
rect 582 482 585 538
rect 582 472 585 478
rect 522 348 526 351
rect 598 351 601 568
rect 614 562 617 568
rect 646 552 649 718
rect 670 702 673 718
rect 710 672 713 678
rect 694 663 697 668
rect 726 662 729 758
rect 734 732 737 747
rect 766 742 769 748
rect 782 741 785 768
rect 810 758 814 761
rect 810 748 814 751
rect 778 738 785 741
rect 802 738 806 741
rect 794 728 798 731
rect 734 672 737 728
rect 782 722 785 728
rect 774 692 777 698
rect 766 662 769 668
rect 646 542 649 548
rect 674 547 678 550
rect 694 491 697 588
rect 726 572 729 658
rect 734 592 737 658
rect 750 552 753 618
rect 758 552 761 568
rect 766 552 769 558
rect 790 552 793 688
rect 822 682 825 868
rect 934 863 937 938
rect 968 903 970 907
rect 974 903 977 907
rect 981 903 984 907
rect 950 872 953 878
rect 862 832 865 858
rect 862 802 865 828
rect 830 762 833 778
rect 862 762 865 778
rect 886 762 889 838
rect 982 812 985 818
rect 830 722 833 728
rect 838 682 841 758
rect 918 752 921 758
rect 982 752 985 808
rect 990 752 993 798
rect 1006 792 1009 818
rect 1030 792 1033 988
rect 1094 952 1097 1148
rect 1102 1132 1105 1148
rect 1102 1063 1105 1118
rect 1102 1052 1105 1059
rect 1118 992 1121 1238
rect 1126 1162 1129 1258
rect 1134 1172 1137 1258
rect 1158 1222 1161 1258
rect 1222 1252 1225 1258
rect 1278 1232 1281 1348
rect 1334 1342 1337 1348
rect 1318 1302 1321 1328
rect 1342 1292 1345 1358
rect 1414 1352 1417 1358
rect 1362 1348 1366 1351
rect 1378 1348 1382 1351
rect 1430 1342 1433 1348
rect 1454 1342 1457 1348
rect 1350 1272 1353 1338
rect 1374 1332 1377 1338
rect 1398 1312 1401 1338
rect 1438 1332 1441 1338
rect 1406 1322 1409 1328
rect 1450 1318 1454 1321
rect 1374 1272 1377 1308
rect 1398 1271 1401 1308
rect 1422 1272 1425 1318
rect 1462 1312 1465 1358
rect 1574 1352 1577 1358
rect 1478 1322 1481 1348
rect 1518 1332 1521 1338
rect 1470 1292 1473 1298
rect 1502 1282 1505 1328
rect 1518 1282 1521 1328
rect 1534 1322 1537 1348
rect 1606 1342 1609 1358
rect 1614 1352 1617 1378
rect 1554 1338 1558 1341
rect 1578 1338 1582 1341
rect 1622 1332 1625 1338
rect 1602 1328 1606 1331
rect 1550 1282 1553 1318
rect 1398 1268 1409 1271
rect 1294 1252 1297 1258
rect 1326 1242 1329 1258
rect 1126 1112 1129 1158
rect 1142 1152 1145 1168
rect 1134 1082 1137 1128
rect 1134 1062 1137 1068
rect 1150 1062 1153 1218
rect 1174 1111 1177 1148
rect 1206 1142 1209 1147
rect 1238 1132 1241 1178
rect 1254 1152 1257 1158
rect 1262 1152 1265 1218
rect 1278 1182 1281 1218
rect 1310 1182 1313 1218
rect 1282 1178 1289 1181
rect 1278 1162 1281 1168
rect 1250 1138 1254 1141
rect 1166 1108 1177 1111
rect 1166 1092 1169 1108
rect 1166 1072 1169 1088
rect 1118 952 1121 978
rect 1078 942 1081 948
rect 1058 928 1062 931
rect 1046 872 1049 918
rect 1070 892 1073 918
rect 1062 872 1065 878
rect 1046 852 1049 859
rect 850 748 854 751
rect 930 748 934 751
rect 858 738 862 741
rect 862 712 865 718
rect 878 692 881 748
rect 886 742 889 748
rect 942 692 945 718
rect 958 702 961 748
rect 966 722 969 748
rect 968 703 970 707
rect 974 703 977 707
rect 981 703 984 707
rect 998 692 1001 788
rect 1030 762 1033 788
rect 1062 771 1065 868
rect 1086 862 1089 948
rect 1094 882 1097 948
rect 1134 942 1137 958
rect 1102 932 1105 938
rect 1150 922 1153 948
rect 1158 942 1161 978
rect 1182 942 1185 988
rect 1194 978 1198 981
rect 1170 938 1174 941
rect 1198 932 1201 938
rect 1110 862 1113 868
rect 1134 862 1137 888
rect 1078 812 1081 818
rect 1062 768 1073 771
rect 978 688 982 691
rect 874 678 878 681
rect 834 659 838 662
rect 886 662 889 688
rect 934 672 937 678
rect 1038 672 1041 678
rect 938 668 942 671
rect 918 663 921 668
rect 874 658 878 661
rect 1054 572 1057 738
rect 1070 682 1073 768
rect 1086 722 1089 858
rect 1110 752 1113 858
rect 1142 792 1145 888
rect 1174 792 1177 878
rect 1190 862 1193 868
rect 1198 852 1201 918
rect 1206 892 1209 958
rect 1214 952 1217 1098
rect 1222 1052 1225 1068
rect 1230 1062 1233 1108
rect 1238 1062 1241 1118
rect 1222 1002 1225 1048
rect 1218 948 1222 951
rect 1230 941 1233 1058
rect 1222 938 1233 941
rect 1214 872 1217 878
rect 1222 862 1225 938
rect 1238 892 1241 1058
rect 1246 932 1249 1088
rect 1262 1062 1265 1108
rect 1286 1072 1289 1178
rect 1310 1162 1313 1168
rect 1350 1152 1353 1268
rect 1366 1262 1369 1268
rect 1382 1252 1385 1258
rect 1394 1248 1398 1251
rect 1406 1212 1409 1268
rect 1430 1262 1433 1268
rect 1438 1262 1441 1268
rect 1502 1262 1505 1278
rect 1458 1258 1462 1261
rect 1306 1148 1310 1151
rect 1294 1142 1297 1148
rect 1358 1142 1361 1158
rect 1374 1152 1377 1158
rect 1354 1138 1358 1141
rect 1306 1058 1310 1061
rect 1254 952 1257 1018
rect 1318 972 1321 1118
rect 1334 1092 1337 1128
rect 1374 1102 1377 1148
rect 1398 1142 1401 1148
rect 1362 1088 1366 1091
rect 1382 1072 1385 1078
rect 1334 952 1337 968
rect 1306 938 1310 941
rect 1254 932 1257 938
rect 1310 922 1313 928
rect 1334 922 1337 938
rect 1282 918 1286 921
rect 1322 918 1326 921
rect 1270 882 1273 888
rect 1238 872 1241 878
rect 1350 872 1353 1068
rect 1414 1062 1417 1258
rect 1430 1192 1433 1208
rect 1422 1132 1425 1148
rect 1438 1111 1441 1258
rect 1478 1252 1481 1258
rect 1454 1212 1457 1248
rect 1480 1203 1482 1207
rect 1486 1203 1489 1207
rect 1493 1203 1496 1207
rect 1502 1172 1505 1218
rect 1518 1152 1521 1278
rect 1526 1262 1529 1268
rect 1550 1262 1553 1268
rect 1558 1242 1561 1248
rect 1566 1242 1569 1318
rect 1590 1291 1593 1318
rect 1590 1288 1601 1291
rect 1590 1272 1593 1278
rect 1574 1262 1577 1268
rect 1574 1242 1577 1258
rect 1586 1248 1590 1251
rect 1430 1108 1441 1111
rect 1422 942 1425 1088
rect 1430 992 1433 1108
rect 1454 1092 1457 1128
rect 1462 1102 1465 1118
rect 1458 1088 1462 1091
rect 1470 1072 1473 1098
rect 1494 1062 1497 1138
rect 1526 1122 1529 1147
rect 1558 1142 1561 1158
rect 1566 1152 1569 1158
rect 1570 1148 1577 1151
rect 1542 1132 1545 1138
rect 1526 1062 1529 1068
rect 1494 1052 1497 1058
rect 1542 1022 1545 1128
rect 1550 1082 1553 1088
rect 1558 1082 1561 1138
rect 1574 1062 1577 1148
rect 1582 1072 1585 1118
rect 1590 1102 1593 1118
rect 1562 1058 1566 1061
rect 1586 1058 1590 1061
rect 1480 1003 1482 1007
rect 1486 1003 1489 1007
rect 1493 1003 1496 1007
rect 1494 951 1497 958
rect 1510 942 1513 1018
rect 1538 988 1542 991
rect 1590 972 1593 1018
rect 1598 952 1601 1288
rect 1606 1252 1609 1268
rect 1630 1262 1633 1268
rect 1618 1258 1622 1261
rect 1638 1252 1641 1358
rect 1758 1352 1761 1468
rect 1810 1428 1814 1431
rect 1830 1352 1833 1468
rect 1918 1462 1921 1548
rect 1846 1452 1849 1459
rect 1906 1428 1910 1431
rect 1910 1372 1913 1378
rect 1650 1348 1654 1351
rect 1690 1348 1694 1351
rect 1662 1342 1665 1348
rect 1842 1348 1846 1351
rect 1726 1342 1729 1347
rect 1658 1338 1662 1341
rect 1674 1338 1678 1341
rect 1646 1332 1649 1338
rect 1662 1272 1665 1338
rect 1670 1322 1673 1328
rect 1686 1292 1689 1338
rect 1670 1272 1673 1278
rect 1606 1082 1609 1248
rect 1638 1192 1641 1248
rect 1654 1222 1657 1258
rect 1718 1252 1721 1268
rect 1758 1262 1761 1348
rect 1830 1342 1833 1348
rect 1778 1258 1782 1261
rect 1686 1162 1689 1168
rect 1650 1147 1654 1150
rect 1646 1122 1649 1147
rect 1670 1132 1673 1138
rect 1622 1082 1625 1098
rect 1626 1078 1630 1081
rect 1606 1062 1609 1078
rect 1646 1072 1649 1088
rect 1670 1072 1673 1078
rect 1618 1068 1622 1071
rect 1674 1068 1678 1071
rect 1686 1062 1689 1068
rect 1634 1058 1638 1061
rect 1658 1058 1662 1061
rect 1662 942 1665 947
rect 1374 882 1377 938
rect 1430 932 1433 938
rect 1394 918 1398 921
rect 1326 862 1329 868
rect 1218 858 1222 861
rect 1258 858 1262 861
rect 1198 822 1201 848
rect 1146 788 1150 791
rect 1190 752 1193 818
rect 1214 762 1217 788
rect 1230 762 1233 858
rect 1214 752 1217 758
rect 1258 748 1262 751
rect 1094 732 1097 748
rect 1110 742 1113 748
rect 1070 663 1073 668
rect 1110 592 1113 718
rect 1166 692 1169 738
rect 1166 682 1169 688
rect 1134 662 1137 678
rect 1190 662 1193 748
rect 1238 672 1241 738
rect 1254 732 1257 738
rect 1270 732 1273 758
rect 1282 738 1286 741
rect 1274 728 1278 731
rect 1226 638 1230 641
rect 1238 632 1241 668
rect 1246 642 1249 718
rect 1334 692 1337 868
rect 1366 742 1369 878
rect 1378 868 1382 871
rect 1390 862 1393 868
rect 1422 862 1425 878
rect 1430 862 1433 908
rect 1454 882 1457 888
rect 1510 872 1513 938
rect 1678 912 1681 1058
rect 1694 952 1697 1128
rect 1718 1112 1721 1238
rect 1726 1162 1729 1218
rect 1718 1062 1721 1108
rect 1734 1092 1737 1148
rect 1742 1142 1745 1238
rect 1774 1172 1777 1258
rect 1790 1252 1793 1318
rect 1750 1151 1753 1168
rect 1790 1152 1793 1218
rect 1798 1152 1801 1158
rect 1742 1082 1745 1138
rect 1766 1132 1769 1138
rect 1806 1132 1809 1338
rect 1894 1331 1897 1348
rect 1894 1328 1902 1331
rect 1886 1282 1889 1288
rect 1842 1278 1846 1281
rect 1870 1261 1873 1278
rect 1918 1272 1921 1348
rect 1866 1258 1873 1261
rect 1890 1258 1894 1261
rect 1914 1258 1918 1261
rect 1830 1242 1833 1258
rect 1862 1182 1865 1258
rect 1866 1178 1873 1181
rect 1822 1152 1825 1178
rect 1830 1152 1833 1158
rect 1838 1152 1841 1158
rect 1862 1152 1865 1158
rect 1850 1148 1854 1151
rect 1846 1138 1854 1141
rect 1806 1092 1809 1128
rect 1846 1092 1849 1138
rect 1854 1132 1857 1138
rect 1726 942 1729 968
rect 1742 952 1745 1078
rect 1750 1052 1753 1068
rect 1870 1062 1873 1178
rect 1878 1162 1881 1168
rect 1894 1152 1897 1238
rect 1902 1152 1905 1258
rect 1926 1242 1929 1248
rect 1934 1242 1937 1278
rect 1886 1142 1889 1148
rect 1894 1142 1897 1148
rect 1894 1092 1897 1138
rect 1906 1128 1910 1131
rect 1918 1102 1921 1148
rect 1942 1092 1945 1618
rect 1950 1542 1953 1548
rect 1950 1342 1953 1348
rect 1950 1262 1953 1268
rect 1918 1082 1921 1088
rect 1902 1062 1905 1068
rect 1826 1058 1830 1061
rect 1806 992 1809 1018
rect 1766 952 1769 958
rect 1502 862 1505 868
rect 1382 852 1385 858
rect 1406 852 1409 858
rect 1374 792 1377 838
rect 1480 803 1482 807
rect 1486 803 1489 807
rect 1493 803 1496 807
rect 1534 792 1537 868
rect 1550 862 1553 908
rect 1598 892 1601 898
rect 1694 882 1697 938
rect 1730 918 1734 921
rect 1694 872 1697 878
rect 1718 872 1721 918
rect 1790 882 1793 948
rect 1838 942 1841 988
rect 1858 947 1862 950
rect 1838 892 1841 938
rect 1914 918 1918 921
rect 1762 878 1766 881
rect 1894 879 1902 881
rect 1894 878 1905 879
rect 1630 868 1638 871
rect 1574 862 1577 868
rect 1586 858 1590 861
rect 1606 852 1609 858
rect 1622 822 1625 868
rect 1630 792 1633 868
rect 1638 842 1641 868
rect 1650 858 1654 861
rect 1662 852 1665 858
rect 1678 852 1681 858
rect 1646 822 1649 828
rect 1654 822 1657 848
rect 1374 782 1377 788
rect 1646 762 1649 818
rect 1662 772 1665 848
rect 1682 838 1686 841
rect 1706 838 1710 841
rect 1734 832 1737 868
rect 1742 862 1745 878
rect 1814 872 1817 878
rect 1754 848 1758 851
rect 1782 832 1785 858
rect 1586 748 1590 751
rect 1650 748 1654 751
rect 1346 738 1350 741
rect 1378 738 1382 741
rect 1398 692 1401 698
rect 1334 682 1337 688
rect 1346 658 1350 661
rect 1406 632 1409 668
rect 1422 662 1425 748
rect 1462 692 1465 738
rect 1478 702 1481 718
rect 834 558 838 561
rect 806 552 809 558
rect 710 542 713 548
rect 726 542 729 548
rect 838 542 841 548
rect 862 542 865 558
rect 870 552 873 558
rect 1038 552 1041 558
rect 1054 552 1057 558
rect 882 548 886 551
rect 1082 548 1086 551
rect 774 532 777 538
rect 878 532 881 538
rect 902 532 905 538
rect 730 528 734 531
rect 842 528 846 531
rect 874 528 878 531
rect 918 528 926 531
rect 710 522 713 528
rect 690 488 697 491
rect 682 478 686 481
rect 638 472 641 478
rect 734 472 737 528
rect 742 462 745 518
rect 786 488 790 491
rect 806 472 809 478
rect 818 468 822 471
rect 830 452 833 478
rect 782 372 785 448
rect 694 352 697 358
rect 510 342 513 348
rect 502 332 505 338
rect 530 328 534 331
rect 542 292 545 338
rect 482 288 486 291
rect 598 281 601 347
rect 678 342 681 348
rect 838 342 841 528
rect 846 442 849 448
rect 854 352 857 518
rect 862 492 865 528
rect 886 492 889 498
rect 902 482 905 528
rect 918 472 921 528
rect 934 492 937 528
rect 878 391 881 468
rect 902 462 905 468
rect 918 452 921 468
rect 926 462 929 468
rect 950 462 953 528
rect 906 448 910 451
rect 878 388 886 391
rect 850 348 854 351
rect 918 351 921 358
rect 722 338 726 341
rect 614 321 617 338
rect 654 322 657 328
rect 614 318 625 321
rect 598 278 609 281
rect 378 258 382 261
rect 510 242 513 268
rect 206 152 209 168
rect 318 152 321 158
rect 350 152 353 168
rect 406 152 409 228
rect 456 203 458 207
rect 462 203 465 207
rect 469 203 472 207
rect 598 192 601 268
rect 606 263 609 278
rect 490 168 494 171
rect 242 148 246 151
rect 334 148 342 151
rect 190 92 193 148
rect 262 132 265 138
rect 270 122 273 148
rect 234 118 238 121
rect 278 111 281 138
rect 286 132 289 138
rect 294 132 297 148
rect 302 122 305 138
rect 270 108 281 111
rect 270 102 273 108
rect 114 68 118 71
rect 178 68 182 71
rect 206 62 209 78
rect 214 72 217 88
rect 270 82 273 98
rect 302 92 305 108
rect 310 92 313 128
rect 334 92 337 148
rect 298 78 302 81
rect 238 72 241 78
rect 310 72 313 88
rect 226 68 230 71
rect 34 58 38 61
rect 154 58 158 61
rect 142 52 145 58
rect 166 52 169 58
rect 50 48 54 51
rect 162 48 166 51
rect 194 48 198 51
rect 254 42 257 58
rect 294 42 297 58
rect 326 52 329 78
rect 342 72 345 128
rect 414 102 417 158
rect 470 152 473 168
rect 430 132 433 138
rect 462 112 465 138
rect 354 88 358 91
rect 414 82 417 98
rect 454 62 457 108
rect 470 92 473 148
rect 550 122 553 148
rect 486 91 489 118
rect 502 92 505 118
rect 486 88 497 91
rect 470 71 473 88
rect 494 82 497 88
rect 466 68 473 71
rect 414 52 417 59
rect 486 52 489 78
rect 518 72 521 78
rect 494 52 497 58
rect 510 52 513 58
rect 534 42 537 58
rect 558 52 561 148
rect 598 142 601 158
rect 594 138 598 141
rect 574 132 577 138
rect 566 79 574 81
rect 606 82 609 88
rect 614 82 617 128
rect 622 102 625 318
rect 662 301 665 328
rect 654 298 665 301
rect 654 262 657 298
rect 678 291 681 328
rect 678 288 686 291
rect 686 282 689 288
rect 694 252 697 278
rect 718 262 721 278
rect 750 262 753 338
rect 786 328 790 331
rect 758 311 761 328
rect 758 308 769 311
rect 766 282 769 308
rect 766 272 769 278
rect 746 258 750 261
rect 770 258 774 261
rect 718 232 721 258
rect 734 242 737 248
rect 782 242 785 328
rect 838 272 841 338
rect 950 332 953 458
rect 958 392 961 538
rect 1030 532 1033 538
rect 978 518 982 521
rect 968 503 970 507
rect 974 503 977 507
rect 981 503 984 507
rect 1002 488 1006 491
rect 990 452 993 458
rect 998 392 1001 478
rect 1014 462 1017 518
rect 1062 482 1065 548
rect 1094 542 1097 548
rect 1066 478 1070 481
rect 1030 462 1033 478
rect 1078 472 1081 528
rect 1074 468 1078 471
rect 978 388 982 391
rect 1018 340 1022 343
rect 1046 342 1049 468
rect 1086 462 1089 538
rect 1102 442 1105 568
rect 1158 562 1161 568
rect 1118 552 1121 558
rect 1138 548 1142 551
rect 1194 548 1201 551
rect 1218 548 1222 551
rect 1126 542 1129 548
rect 1174 542 1177 548
rect 1198 542 1201 548
rect 1294 542 1297 618
rect 1398 582 1401 618
rect 1470 592 1473 658
rect 1502 642 1505 748
rect 1550 732 1553 738
rect 1630 732 1633 738
rect 1526 722 1529 728
rect 1550 692 1553 728
rect 1638 712 1641 748
rect 1662 742 1665 758
rect 1670 742 1673 818
rect 1682 758 1686 761
rect 1702 752 1705 758
rect 1718 738 1726 741
rect 1638 692 1641 708
rect 1606 672 1609 678
rect 1646 672 1649 738
rect 1690 728 1694 731
rect 1654 722 1657 728
rect 1674 718 1678 721
rect 1662 672 1665 688
rect 1718 682 1721 738
rect 1694 672 1697 678
rect 1546 668 1550 671
rect 1626 668 1630 671
rect 1590 662 1593 668
rect 1538 658 1542 661
rect 1546 658 1550 661
rect 1598 642 1601 668
rect 1646 662 1649 668
rect 1646 652 1649 658
rect 1480 603 1482 607
rect 1486 603 1489 607
rect 1493 603 1496 607
rect 1302 542 1305 548
rect 1134 538 1142 541
rect 1210 538 1214 541
rect 1134 532 1137 538
rect 1182 532 1185 538
rect 1118 492 1121 508
rect 1134 472 1137 528
rect 1062 352 1065 388
rect 1102 352 1105 438
rect 1034 338 1038 341
rect 918 272 921 328
rect 968 303 970 307
rect 974 303 977 307
rect 981 303 984 307
rect 958 272 961 278
rect 990 272 993 338
rect 1042 328 1046 331
rect 1054 322 1057 338
rect 1118 332 1121 368
rect 1126 332 1129 368
rect 1134 342 1137 468
rect 1142 362 1145 518
rect 1150 492 1153 528
rect 1190 521 1193 538
rect 1182 518 1193 521
rect 1182 492 1185 518
rect 1190 482 1193 488
rect 1198 472 1201 488
rect 1154 458 1158 461
rect 1158 452 1161 458
rect 1086 282 1089 308
rect 1054 272 1057 278
rect 754 238 758 241
rect 742 232 745 238
rect 786 218 790 221
rect 758 172 761 178
rect 670 142 673 158
rect 694 152 697 168
rect 778 158 782 161
rect 650 138 654 141
rect 638 92 641 108
rect 566 78 577 79
rect 566 62 569 78
rect 618 68 622 71
rect 590 62 593 68
rect 598 62 601 68
rect 638 52 641 58
rect 546 48 550 51
rect 456 3 458 7
rect 462 3 465 7
rect 469 3 472 7
rect 574 -19 578 -18
rect 582 -19 585 18
rect 574 -22 585 -19
rect 654 -18 657 138
rect 670 82 673 98
rect 694 62 697 148
rect 750 122 753 158
rect 742 118 750 121
rect 742 82 745 118
rect 774 92 777 148
rect 806 142 809 218
rect 814 192 817 238
rect 846 192 849 259
rect 874 218 878 221
rect 918 192 921 218
rect 934 192 937 258
rect 1022 212 1025 218
rect 1086 202 1089 259
rect 878 182 881 188
rect 814 152 817 158
rect 886 152 889 158
rect 810 138 814 141
rect 750 82 753 88
rect 782 82 785 128
rect 790 122 793 138
rect 838 132 841 138
rect 826 128 830 131
rect 798 112 801 128
rect 814 102 817 118
rect 822 112 825 118
rect 814 92 817 98
rect 790 82 793 88
rect 822 82 825 108
rect 862 102 865 138
rect 870 92 873 138
rect 902 122 905 148
rect 918 142 921 148
rect 914 138 918 141
rect 930 128 934 131
rect 942 131 945 148
rect 1006 142 1009 148
rect 942 128 950 131
rect 990 122 993 138
rect 1006 122 1009 128
rect 968 103 970 107
rect 974 103 977 107
rect 981 103 984 107
rect 866 88 870 91
rect 918 82 921 88
rect 790 72 793 78
rect 798 72 801 78
rect 770 68 774 71
rect 882 68 886 71
rect 854 62 857 68
rect 926 62 929 78
rect 998 72 1001 118
rect 1038 112 1041 138
rect 1050 118 1054 121
rect 1062 112 1065 158
rect 1094 152 1097 158
rect 1102 152 1105 328
rect 1182 282 1185 368
rect 1190 351 1193 358
rect 1206 352 1209 538
rect 1214 442 1217 528
rect 1242 518 1246 521
rect 1278 472 1281 538
rect 1366 532 1369 548
rect 1350 472 1353 518
rect 1374 492 1377 528
rect 1390 512 1393 538
rect 1406 532 1409 578
rect 1394 488 1398 491
rect 1438 482 1441 558
rect 1450 548 1454 551
rect 1470 542 1473 548
rect 1478 532 1481 568
rect 1494 562 1497 578
rect 1510 491 1513 548
rect 1526 542 1529 548
rect 1590 542 1593 548
rect 1502 488 1513 491
rect 1518 532 1521 538
rect 1502 482 1505 488
rect 1510 472 1513 478
rect 1214 372 1217 438
rect 1246 392 1249 468
rect 1262 463 1265 468
rect 1238 352 1241 358
rect 1302 352 1305 468
rect 1330 458 1334 461
rect 1446 392 1449 468
rect 1454 463 1457 468
rect 1518 462 1521 528
rect 1526 492 1529 538
rect 1558 532 1562 535
rect 1566 522 1569 532
rect 1530 478 1534 481
rect 1526 462 1529 468
rect 1558 462 1561 518
rect 1566 492 1569 518
rect 1598 512 1601 638
rect 1606 632 1609 648
rect 1634 638 1638 641
rect 1622 592 1625 628
rect 1630 562 1633 568
rect 1606 552 1609 558
rect 1638 552 1641 578
rect 1614 532 1617 538
rect 1586 488 1590 491
rect 1582 462 1585 488
rect 1546 458 1550 461
rect 1570 458 1574 461
rect 1562 438 1566 441
rect 1480 403 1482 407
rect 1486 403 1489 407
rect 1493 403 1496 407
rect 1354 368 1361 371
rect 1358 352 1361 368
rect 1514 348 1518 351
rect 1390 342 1393 348
rect 1206 312 1209 338
rect 1222 292 1225 328
rect 1294 312 1297 338
rect 1238 292 1241 308
rect 1350 272 1353 308
rect 1390 272 1393 338
rect 1446 322 1449 338
rect 1446 272 1449 318
rect 1290 268 1294 271
rect 1490 258 1494 261
rect 1118 212 1121 218
rect 1110 192 1113 198
rect 1074 138 1078 141
rect 1118 132 1121 208
rect 1054 92 1057 108
rect 1034 88 1038 91
rect 1006 82 1009 88
rect 1118 72 1121 128
rect 1134 72 1137 238
rect 1174 202 1177 258
rect 1334 252 1337 258
rect 1374 242 1377 258
rect 1238 191 1241 218
rect 1238 188 1249 191
rect 1246 152 1249 188
rect 1338 158 1342 161
rect 1394 158 1398 161
rect 1178 148 1185 151
rect 1150 112 1153 148
rect 1158 102 1161 118
rect 1182 92 1185 148
rect 1278 151 1281 158
rect 1190 142 1193 148
rect 1206 102 1209 118
rect 1010 68 1014 71
rect 1022 62 1025 68
rect 1046 62 1049 68
rect 1070 62 1073 68
rect 1150 63 1153 78
rect 1198 62 1201 68
rect 1206 62 1209 98
rect 1230 92 1233 128
rect 1214 82 1217 88
rect 1226 78 1230 81
rect 1246 72 1249 78
rect 874 48 878 51
rect 854 42 857 48
rect 982 42 985 58
rect 1030 42 1033 48
rect 1070 42 1073 58
rect 1086 42 1089 58
rect 1182 52 1185 58
rect 1222 52 1225 68
rect 1230 52 1233 58
rect 1254 52 1257 148
rect 1310 132 1313 138
rect 1318 122 1321 148
rect 1262 72 1265 88
rect 1294 72 1297 78
rect 1318 62 1321 118
rect 1266 58 1270 61
rect 1278 52 1281 58
rect 1334 52 1337 158
rect 1414 152 1417 238
rect 1430 192 1433 218
rect 1454 151 1457 238
rect 1486 222 1489 258
rect 1480 203 1482 207
rect 1486 203 1489 207
rect 1493 203 1496 207
rect 1502 172 1505 328
rect 1550 292 1553 428
rect 1566 392 1569 438
rect 1574 432 1577 448
rect 1614 442 1617 528
rect 1582 332 1585 338
rect 1546 288 1550 291
rect 1574 252 1577 259
rect 1522 188 1526 191
rect 1350 102 1353 148
rect 1366 142 1369 148
rect 1358 122 1361 138
rect 1374 102 1377 148
rect 1390 142 1393 148
rect 1398 112 1401 148
rect 1406 122 1409 138
rect 1422 132 1425 138
rect 1370 88 1374 91
rect 1390 62 1393 98
rect 1398 91 1401 108
rect 1414 92 1417 118
rect 1398 88 1406 91
rect 1438 82 1441 148
rect 1542 142 1545 158
rect 1554 148 1558 151
rect 1582 142 1585 328
rect 1598 262 1601 438
rect 1622 352 1625 498
rect 1646 492 1649 548
rect 1654 522 1657 538
rect 1662 472 1665 668
rect 1702 662 1705 668
rect 1694 642 1697 648
rect 1670 582 1673 618
rect 1702 562 1705 578
rect 1710 562 1713 578
rect 1718 572 1721 628
rect 1718 562 1721 568
rect 1670 552 1673 558
rect 1694 552 1697 558
rect 1710 542 1713 548
rect 1726 542 1729 738
rect 1734 732 1737 768
rect 1742 752 1745 818
rect 1782 772 1785 818
rect 1762 728 1766 731
rect 1734 702 1737 728
rect 1734 682 1737 698
rect 1758 671 1761 718
rect 1774 712 1777 728
rect 1758 668 1766 671
rect 1782 662 1785 718
rect 1790 692 1793 858
rect 1806 762 1809 768
rect 1798 752 1801 758
rect 1838 732 1841 848
rect 1862 832 1865 868
rect 1894 862 1897 878
rect 1918 862 1921 908
rect 1926 902 1929 948
rect 1942 942 1945 948
rect 1950 912 1953 1218
rect 1946 868 1950 871
rect 1886 841 1889 858
rect 1882 838 1889 841
rect 1854 742 1857 748
rect 1838 692 1841 728
rect 1790 682 1793 688
rect 1806 672 1809 678
rect 1870 672 1873 747
rect 1882 688 1886 691
rect 1822 663 1825 668
rect 1738 658 1742 661
rect 1754 658 1758 661
rect 1738 648 1742 651
rect 1766 651 1769 658
rect 1762 648 1769 651
rect 1894 641 1897 658
rect 1910 642 1913 648
rect 1894 638 1902 641
rect 1782 572 1785 618
rect 1802 558 1806 561
rect 1754 548 1758 551
rect 1770 548 1774 551
rect 1862 551 1865 568
rect 1770 538 1774 541
rect 1786 538 1790 541
rect 1642 459 1646 462
rect 1678 452 1681 538
rect 1730 528 1734 531
rect 1686 502 1689 518
rect 1690 478 1694 481
rect 1698 478 1702 481
rect 1690 468 1694 471
rect 1718 462 1721 498
rect 1706 458 1710 461
rect 1682 448 1686 451
rect 1662 392 1665 438
rect 1734 352 1737 468
rect 1750 463 1753 468
rect 1782 432 1785 528
rect 1798 462 1801 548
rect 1822 542 1825 548
rect 1870 542 1873 638
rect 1918 602 1921 658
rect 1926 592 1929 698
rect 1934 692 1937 718
rect 1946 668 1950 671
rect 1934 592 1937 598
rect 1806 502 1809 518
rect 1810 488 1814 491
rect 1682 348 1686 351
rect 1754 348 1758 351
rect 1734 342 1737 348
rect 1670 292 1673 328
rect 1678 292 1681 298
rect 1650 288 1654 291
rect 1622 282 1625 288
rect 1686 282 1689 338
rect 1702 302 1705 318
rect 1670 272 1673 278
rect 1546 138 1550 141
rect 1546 128 1550 131
rect 1446 62 1449 88
rect 1454 82 1457 128
rect 1502 92 1505 98
rect 1574 62 1577 138
rect 1582 122 1585 128
rect 1598 101 1601 258
rect 1590 98 1601 101
rect 1582 62 1585 88
rect 1590 82 1593 98
rect 1622 92 1625 118
rect 1622 82 1625 88
rect 1630 82 1633 148
rect 1646 142 1649 248
rect 1686 162 1689 268
rect 1742 263 1745 348
rect 1822 292 1825 347
rect 1786 288 1790 291
rect 1774 282 1777 288
rect 1714 258 1718 261
rect 1774 192 1777 278
rect 1806 262 1809 268
rect 1822 263 1825 288
rect 1822 258 1825 259
rect 1738 188 1742 191
rect 1762 158 1766 161
rect 1686 152 1689 158
rect 1730 148 1734 151
rect 1674 118 1678 121
rect 1646 79 1654 81
rect 1646 78 1657 79
rect 1590 72 1593 78
rect 1646 62 1649 78
rect 1670 72 1673 88
rect 1634 58 1638 61
rect 1674 58 1678 61
rect 1686 61 1689 118
rect 1682 58 1689 61
rect 1694 52 1697 138
rect 1702 122 1705 138
rect 1710 61 1713 148
rect 1782 142 1785 158
rect 1790 152 1793 258
rect 1830 251 1833 538
rect 1938 528 1942 531
rect 1910 492 1913 528
rect 1854 462 1857 468
rect 1918 462 1921 508
rect 1822 248 1833 251
rect 1798 152 1801 158
rect 1774 122 1777 138
rect 1806 122 1809 138
rect 1814 132 1817 148
rect 1726 92 1729 118
rect 1758 92 1761 118
rect 1822 82 1825 248
rect 1846 192 1849 458
rect 1870 372 1873 458
rect 1894 368 1902 371
rect 1870 191 1873 368
rect 1894 352 1897 368
rect 1918 331 1921 348
rect 1918 328 1926 331
rect 1886 292 1889 318
rect 1906 279 1913 281
rect 1902 278 1913 279
rect 1910 262 1913 278
rect 1918 241 1921 258
rect 1918 238 1926 241
rect 1862 188 1873 191
rect 1834 148 1838 151
rect 1862 142 1865 188
rect 1886 162 1889 218
rect 1838 132 1841 138
rect 1830 122 1833 128
rect 1838 82 1841 128
rect 1718 72 1721 78
rect 1758 62 1761 68
rect 1782 62 1785 78
rect 1854 72 1857 78
rect 1878 62 1881 147
rect 1942 122 1945 128
rect 1942 92 1945 118
rect 1710 58 1718 61
rect 1822 52 1825 58
rect 1258 48 1262 51
rect 1630 42 1633 48
rect 846 32 849 38
rect 766 -18 769 18
rect 1480 3 1482 7
rect 1486 3 1489 7
rect 1493 3 1496 7
rect 654 -22 658 -18
rect 766 -22 770 -18
<< m3contact >>
rect 970 1703 974 1707
rect 977 1703 981 1707
rect 1062 1698 1066 1702
rect 1078 1688 1082 1692
rect 6 1678 10 1682
rect 62 1678 66 1682
rect 94 1678 98 1682
rect 126 1678 130 1682
rect 134 1678 138 1682
rect 206 1678 210 1682
rect 214 1678 218 1682
rect 406 1678 410 1682
rect 430 1678 434 1682
rect 622 1678 626 1682
rect 1062 1678 1066 1682
rect 22 1668 26 1672
rect 54 1658 58 1662
rect 30 1648 34 1652
rect 110 1668 114 1672
rect 86 1658 90 1662
rect 118 1658 122 1662
rect 70 1638 74 1642
rect 102 1638 106 1642
rect 182 1668 186 1672
rect 166 1658 170 1662
rect 150 1648 154 1652
rect 142 1638 146 1642
rect 62 1468 66 1472
rect 14 1438 18 1442
rect 70 1398 74 1402
rect 6 1358 10 1362
rect 62 1338 66 1342
rect 62 1298 66 1302
rect 14 1238 18 1242
rect 294 1648 298 1652
rect 262 1638 266 1642
rect 238 1618 242 1622
rect 254 1618 258 1622
rect 390 1648 394 1652
rect 318 1618 322 1622
rect 358 1558 362 1562
rect 374 1558 378 1562
rect 166 1548 170 1552
rect 198 1548 202 1552
rect 142 1538 146 1542
rect 110 1468 114 1472
rect 118 1468 122 1472
rect 142 1458 146 1462
rect 86 1278 90 1282
rect 134 1438 138 1442
rect 190 1538 194 1542
rect 238 1538 242 1542
rect 206 1508 210 1512
rect 238 1478 242 1482
rect 414 1551 418 1552
rect 414 1548 418 1551
rect 286 1538 290 1542
rect 302 1518 306 1522
rect 310 1498 314 1502
rect 254 1458 258 1462
rect 182 1418 186 1422
rect 158 1368 162 1372
rect 126 1348 130 1352
rect 134 1338 138 1342
rect 142 1328 146 1332
rect 142 1268 146 1272
rect 190 1358 194 1362
rect 198 1338 202 1342
rect 254 1398 258 1402
rect 230 1358 234 1362
rect 222 1338 226 1342
rect 190 1328 194 1332
rect 206 1328 210 1332
rect 214 1328 218 1332
rect 166 1268 170 1272
rect 158 1258 162 1262
rect 86 1238 90 1242
rect 102 1168 106 1172
rect 126 1148 130 1152
rect 134 1148 138 1152
rect 102 1138 106 1142
rect 118 1138 122 1142
rect 142 1140 146 1144
rect 190 1128 194 1132
rect 110 1088 114 1092
rect 158 1088 162 1092
rect 78 1078 82 1082
rect 86 1078 90 1082
rect 126 1078 130 1082
rect 150 1078 154 1082
rect 14 1068 18 1072
rect 78 1068 82 1072
rect 22 1038 26 1042
rect 54 1038 58 1042
rect 14 958 18 962
rect 22 958 26 962
rect 6 948 10 952
rect 22 948 26 952
rect 38 908 42 912
rect 22 898 26 902
rect 14 868 18 872
rect 110 1068 114 1072
rect 166 1078 170 1082
rect 174 1078 178 1082
rect 102 1058 106 1062
rect 134 1058 138 1062
rect 126 1048 130 1052
rect 142 1048 146 1052
rect 150 1018 154 1022
rect 142 988 146 992
rect 78 938 82 942
rect 54 898 58 902
rect 78 928 82 932
rect 126 928 130 932
rect 86 918 90 922
rect 102 918 106 922
rect 62 868 66 872
rect 118 908 122 912
rect 134 898 138 902
rect 78 848 82 852
rect 102 798 106 802
rect 118 798 122 802
rect 62 788 66 792
rect 94 788 98 792
rect 6 748 10 752
rect 54 748 58 752
rect 70 748 74 752
rect 94 748 98 752
rect 30 738 34 742
rect 70 738 74 742
rect 94 728 98 732
rect 6 648 10 652
rect 30 628 34 632
rect 14 538 18 542
rect 30 538 34 542
rect 94 568 98 572
rect 102 558 106 562
rect 110 538 114 542
rect 38 488 42 492
rect 6 448 10 452
rect 14 388 18 392
rect 86 478 90 482
rect 70 358 74 362
rect 110 488 114 492
rect 126 558 130 562
rect 246 1328 250 1332
rect 238 1318 242 1322
rect 270 1418 274 1422
rect 286 1398 290 1402
rect 270 1358 274 1362
rect 302 1348 306 1352
rect 430 1668 434 1672
rect 438 1668 442 1672
rect 574 1668 578 1672
rect 622 1668 626 1672
rect 694 1668 698 1672
rect 478 1658 482 1662
rect 614 1658 618 1662
rect 662 1658 666 1662
rect 494 1648 498 1652
rect 470 1618 474 1622
rect 518 1618 522 1622
rect 458 1603 462 1607
rect 465 1603 469 1607
rect 446 1578 450 1582
rect 606 1638 610 1642
rect 646 1638 650 1642
rect 630 1618 634 1622
rect 566 1588 570 1592
rect 550 1558 554 1562
rect 510 1538 514 1542
rect 430 1518 434 1522
rect 470 1518 474 1522
rect 422 1498 426 1502
rect 334 1478 338 1482
rect 526 1518 530 1522
rect 598 1528 602 1532
rect 582 1518 586 1522
rect 606 1518 610 1522
rect 566 1508 570 1512
rect 574 1508 578 1512
rect 510 1498 514 1502
rect 534 1488 538 1492
rect 366 1468 370 1472
rect 398 1468 402 1472
rect 422 1468 426 1472
rect 438 1468 442 1472
rect 518 1468 522 1472
rect 374 1458 378 1462
rect 374 1448 378 1452
rect 358 1388 362 1392
rect 414 1458 418 1462
rect 390 1438 394 1442
rect 422 1438 426 1442
rect 382 1428 386 1432
rect 382 1368 386 1372
rect 318 1348 322 1352
rect 326 1338 330 1342
rect 302 1328 306 1332
rect 350 1338 354 1342
rect 286 1308 290 1312
rect 342 1308 346 1312
rect 302 1278 306 1282
rect 342 1278 346 1282
rect 294 1268 298 1272
rect 302 1268 306 1272
rect 334 1268 338 1272
rect 238 1258 242 1262
rect 334 1258 338 1262
rect 334 1238 338 1242
rect 286 1168 290 1172
rect 286 1158 290 1162
rect 614 1508 618 1512
rect 630 1478 634 1482
rect 446 1458 450 1462
rect 510 1458 514 1462
rect 526 1458 530 1462
rect 574 1458 578 1462
rect 458 1403 462 1407
rect 465 1403 469 1407
rect 558 1448 562 1452
rect 518 1438 522 1442
rect 518 1398 522 1402
rect 542 1398 546 1402
rect 574 1398 578 1402
rect 438 1358 442 1362
rect 422 1338 426 1342
rect 374 1328 378 1332
rect 390 1328 394 1332
rect 374 1308 378 1312
rect 438 1338 442 1342
rect 430 1308 434 1312
rect 406 1298 410 1302
rect 430 1288 434 1292
rect 422 1278 426 1282
rect 382 1268 386 1272
rect 374 1248 378 1252
rect 254 1148 258 1152
rect 350 1148 354 1152
rect 358 1138 362 1142
rect 318 1128 322 1132
rect 254 1108 258 1112
rect 238 1088 242 1092
rect 294 1078 298 1082
rect 238 1068 242 1072
rect 302 1058 306 1062
rect 318 1058 322 1062
rect 350 1058 354 1062
rect 198 1048 202 1052
rect 222 1048 226 1052
rect 190 1038 194 1042
rect 262 1018 266 1022
rect 190 947 194 951
rect 150 818 154 822
rect 166 818 170 822
rect 166 748 170 752
rect 142 738 146 742
rect 318 978 322 982
rect 278 948 282 952
rect 310 948 314 952
rect 262 938 266 942
rect 302 928 306 932
rect 270 918 274 922
rect 366 1088 370 1092
rect 438 1268 442 1272
rect 566 1358 570 1362
rect 558 1338 562 1342
rect 478 1288 482 1292
rect 486 1288 490 1292
rect 526 1318 530 1322
rect 542 1318 546 1322
rect 510 1298 514 1302
rect 518 1288 522 1292
rect 526 1268 530 1272
rect 526 1258 530 1262
rect 398 1248 402 1252
rect 422 1248 426 1252
rect 390 1238 394 1242
rect 406 1238 410 1242
rect 502 1248 506 1252
rect 458 1203 462 1207
rect 465 1203 469 1207
rect 478 1198 482 1202
rect 398 1178 402 1182
rect 422 1168 426 1172
rect 438 1168 442 1172
rect 486 1168 490 1172
rect 518 1188 522 1192
rect 518 1168 522 1172
rect 566 1308 570 1312
rect 558 1258 562 1262
rect 558 1248 562 1252
rect 550 1208 554 1212
rect 574 1298 578 1302
rect 590 1458 594 1462
rect 726 1648 730 1652
rect 726 1558 730 1562
rect 694 1528 698 1532
rect 670 1508 674 1512
rect 710 1508 714 1512
rect 686 1498 690 1502
rect 710 1488 714 1492
rect 670 1468 674 1472
rect 630 1438 634 1442
rect 638 1428 642 1432
rect 662 1408 666 1412
rect 774 1538 778 1542
rect 774 1528 778 1532
rect 782 1468 786 1472
rect 630 1388 634 1392
rect 718 1448 722 1452
rect 734 1428 738 1432
rect 750 1418 754 1422
rect 806 1628 810 1632
rect 822 1628 826 1632
rect 870 1658 874 1662
rect 894 1658 898 1662
rect 870 1551 874 1552
rect 870 1548 874 1551
rect 846 1538 850 1542
rect 806 1508 810 1512
rect 822 1478 826 1482
rect 846 1478 850 1482
rect 974 1668 978 1672
rect 1006 1658 1010 1662
rect 1022 1648 1026 1652
rect 1038 1648 1042 1652
rect 942 1628 946 1632
rect 918 1618 922 1622
rect 1078 1618 1082 1622
rect 1158 1698 1162 1702
rect 1326 1698 1330 1702
rect 1510 1698 1514 1702
rect 1526 1698 1530 1702
rect 1150 1678 1154 1682
rect 1382 1678 1386 1682
rect 1446 1678 1450 1682
rect 1270 1668 1274 1672
rect 1390 1668 1394 1672
rect 1454 1668 1458 1672
rect 1470 1668 1474 1672
rect 1510 1668 1514 1672
rect 1118 1658 1122 1662
rect 1150 1658 1154 1662
rect 1118 1648 1122 1652
rect 1110 1618 1114 1622
rect 1070 1608 1074 1612
rect 990 1568 994 1572
rect 1030 1568 1034 1572
rect 910 1558 914 1562
rect 950 1558 954 1562
rect 1014 1558 1018 1562
rect 1246 1628 1250 1632
rect 1318 1628 1322 1632
rect 1190 1598 1194 1602
rect 1270 1598 1274 1602
rect 1294 1598 1298 1602
rect 1214 1578 1218 1582
rect 1182 1558 1186 1562
rect 1238 1558 1242 1562
rect 1286 1558 1290 1562
rect 1310 1578 1314 1582
rect 958 1548 962 1552
rect 998 1548 1002 1552
rect 1022 1548 1026 1552
rect 1086 1548 1090 1552
rect 1150 1548 1154 1552
rect 1214 1548 1218 1552
rect 1262 1548 1266 1552
rect 1278 1548 1282 1552
rect 926 1538 930 1542
rect 902 1528 906 1532
rect 910 1488 914 1492
rect 862 1468 866 1472
rect 886 1468 890 1472
rect 798 1459 802 1463
rect 966 1528 970 1532
rect 1014 1528 1018 1532
rect 1038 1528 1042 1532
rect 1086 1528 1090 1532
rect 970 1503 974 1507
rect 977 1503 981 1507
rect 1046 1488 1050 1492
rect 1030 1478 1034 1482
rect 1038 1478 1042 1482
rect 838 1458 842 1462
rect 870 1458 874 1462
rect 918 1458 922 1462
rect 942 1458 946 1462
rect 966 1458 970 1462
rect 990 1458 994 1462
rect 806 1438 810 1442
rect 830 1438 834 1442
rect 854 1438 858 1442
rect 702 1378 706 1382
rect 662 1368 666 1372
rect 614 1358 618 1362
rect 638 1358 642 1362
rect 630 1348 634 1352
rect 590 1338 594 1342
rect 614 1338 618 1342
rect 598 1278 602 1282
rect 566 1198 570 1202
rect 454 1158 458 1162
rect 502 1158 506 1162
rect 550 1158 554 1162
rect 494 1148 498 1152
rect 406 1138 410 1142
rect 390 1118 394 1122
rect 382 1098 386 1102
rect 398 1098 402 1102
rect 374 1078 378 1082
rect 366 1068 370 1072
rect 350 968 354 972
rect 358 968 362 972
rect 334 958 338 962
rect 406 1078 410 1082
rect 542 1148 546 1152
rect 510 1138 514 1142
rect 654 1338 658 1342
rect 654 1318 658 1322
rect 638 1308 642 1312
rect 678 1348 682 1352
rect 710 1368 714 1372
rect 718 1368 722 1372
rect 742 1368 746 1372
rect 814 1418 818 1422
rect 886 1448 890 1452
rect 862 1428 866 1432
rect 902 1428 906 1432
rect 902 1408 906 1412
rect 694 1348 698 1352
rect 710 1348 714 1352
rect 846 1348 850 1352
rect 726 1338 730 1342
rect 734 1338 738 1342
rect 686 1318 690 1322
rect 630 1258 634 1262
rect 590 1238 594 1242
rect 598 1158 602 1162
rect 622 1158 626 1162
rect 582 1148 586 1152
rect 614 1148 618 1152
rect 566 1128 570 1132
rect 574 1118 578 1122
rect 510 1108 514 1112
rect 414 1068 418 1072
rect 430 1068 434 1072
rect 406 1048 410 1052
rect 390 1038 394 1042
rect 422 1038 426 1042
rect 398 988 402 992
rect 382 958 386 962
rect 374 948 378 952
rect 390 948 394 952
rect 334 938 338 942
rect 358 938 362 942
rect 342 928 346 932
rect 342 918 346 922
rect 270 908 274 912
rect 318 908 322 912
rect 550 1068 554 1072
rect 478 1058 482 1062
rect 462 1038 466 1042
rect 534 1018 538 1022
rect 458 1003 462 1007
rect 465 1003 469 1007
rect 446 968 450 972
rect 542 1008 546 1012
rect 542 978 546 982
rect 534 968 538 972
rect 470 948 474 952
rect 518 948 522 952
rect 382 938 386 942
rect 398 938 402 942
rect 414 938 418 942
rect 390 928 394 932
rect 366 898 370 902
rect 566 978 570 982
rect 558 958 562 962
rect 430 938 434 942
rect 478 938 482 942
rect 430 928 434 932
rect 462 928 466 932
rect 422 918 426 922
rect 406 898 410 902
rect 326 878 330 882
rect 350 878 354 882
rect 382 878 386 882
rect 238 868 242 872
rect 286 868 290 872
rect 230 718 234 722
rect 302 858 306 862
rect 254 828 258 832
rect 182 658 186 662
rect 158 648 162 652
rect 198 638 202 642
rect 182 618 186 622
rect 222 618 226 622
rect 286 818 290 822
rect 358 868 362 872
rect 358 848 362 852
rect 334 818 338 822
rect 318 768 322 772
rect 310 758 314 762
rect 286 728 290 732
rect 302 718 306 722
rect 270 668 274 672
rect 198 568 202 572
rect 254 568 258 572
rect 230 558 234 562
rect 142 538 146 542
rect 222 538 226 542
rect 246 538 250 542
rect 238 528 242 532
rect 182 498 186 502
rect 134 478 138 482
rect 158 478 162 482
rect 214 498 218 502
rect 286 648 290 652
rect 278 638 282 642
rect 294 618 298 622
rect 342 808 346 812
rect 374 848 378 852
rect 446 888 450 892
rect 438 878 442 882
rect 454 878 458 882
rect 446 868 450 872
rect 486 918 490 922
rect 558 918 562 922
rect 518 898 522 902
rect 534 878 538 882
rect 478 868 482 872
rect 422 858 426 862
rect 470 858 474 862
rect 430 848 434 852
rect 462 848 466 852
rect 414 838 418 842
rect 422 808 426 812
rect 458 803 462 807
rect 465 803 469 807
rect 390 788 394 792
rect 454 768 458 772
rect 430 758 434 762
rect 630 1138 634 1142
rect 606 1128 610 1132
rect 710 1328 714 1332
rect 750 1328 754 1332
rect 670 1258 674 1262
rect 694 1258 698 1262
rect 678 1248 682 1252
rect 670 1228 674 1232
rect 694 1228 698 1232
rect 654 1168 658 1172
rect 686 1168 690 1172
rect 718 1318 722 1322
rect 726 1288 730 1292
rect 718 1278 722 1282
rect 726 1248 730 1252
rect 798 1268 802 1272
rect 782 1238 786 1242
rect 798 1238 802 1242
rect 766 1228 770 1232
rect 758 1178 762 1182
rect 710 1148 714 1152
rect 798 1168 802 1172
rect 854 1338 858 1342
rect 838 1318 842 1322
rect 838 1298 842 1302
rect 830 1288 834 1292
rect 838 1278 842 1282
rect 830 1248 834 1252
rect 814 1198 818 1202
rect 878 1308 882 1312
rect 886 1308 890 1312
rect 854 1258 858 1262
rect 870 1258 874 1262
rect 886 1248 890 1252
rect 870 1178 874 1182
rect 838 1168 842 1172
rect 806 1158 810 1162
rect 862 1158 866 1162
rect 838 1148 842 1152
rect 814 1138 818 1142
rect 774 1128 778 1132
rect 622 1108 626 1112
rect 614 1078 618 1082
rect 590 1058 594 1062
rect 598 1048 602 1052
rect 606 1038 610 1042
rect 606 978 610 982
rect 582 948 586 952
rect 598 948 602 952
rect 622 948 626 952
rect 662 1118 666 1122
rect 670 1118 674 1122
rect 678 1108 682 1112
rect 662 1088 666 1092
rect 638 1078 642 1082
rect 646 1078 650 1082
rect 654 1068 658 1072
rect 670 1068 674 1072
rect 766 1098 770 1102
rect 822 1088 826 1092
rect 862 1138 866 1142
rect 854 1118 858 1122
rect 894 1108 898 1112
rect 942 1448 946 1452
rect 934 1428 938 1432
rect 934 1348 938 1352
rect 966 1348 970 1352
rect 918 1338 922 1342
rect 970 1303 974 1307
rect 977 1303 981 1307
rect 1006 1378 1010 1382
rect 1014 1358 1018 1362
rect 958 1258 962 1262
rect 910 1238 914 1242
rect 910 1128 914 1132
rect 934 1128 938 1132
rect 982 1128 986 1132
rect 870 1098 874 1102
rect 902 1098 906 1102
rect 870 1088 874 1092
rect 894 1088 898 1092
rect 702 1078 706 1082
rect 774 1078 778 1082
rect 646 1058 650 1062
rect 662 1058 666 1062
rect 678 1058 682 1062
rect 686 1058 690 1062
rect 750 1058 754 1062
rect 702 1048 706 1052
rect 734 1038 738 1042
rect 774 1028 778 1032
rect 734 1008 738 1012
rect 734 958 738 962
rect 678 948 682 952
rect 686 938 690 942
rect 590 928 594 932
rect 614 928 618 932
rect 630 928 634 932
rect 582 908 586 912
rect 574 898 578 902
rect 582 888 586 892
rect 630 888 634 892
rect 678 888 682 892
rect 686 868 690 872
rect 606 858 610 862
rect 662 858 666 862
rect 590 838 594 842
rect 486 768 490 772
rect 558 768 562 772
rect 374 747 378 751
rect 422 748 426 752
rect 478 748 482 752
rect 366 738 370 742
rect 398 728 402 732
rect 382 698 386 702
rect 374 668 378 672
rect 334 648 338 652
rect 366 618 370 622
rect 350 598 354 602
rect 318 558 322 562
rect 430 738 434 742
rect 478 728 482 732
rect 422 708 426 712
rect 510 758 514 762
rect 534 758 538 762
rect 566 748 570 752
rect 598 748 602 752
rect 558 738 562 742
rect 574 738 578 742
rect 654 768 658 772
rect 630 738 634 742
rect 502 728 506 732
rect 518 728 522 732
rect 534 728 538 732
rect 574 728 578 732
rect 598 728 602 732
rect 534 698 538 702
rect 526 678 530 682
rect 550 678 554 682
rect 542 668 546 672
rect 414 658 418 662
rect 430 658 434 662
rect 502 658 506 662
rect 566 658 570 662
rect 382 598 386 602
rect 358 558 362 562
rect 374 558 378 562
rect 398 558 402 562
rect 622 708 626 712
rect 630 698 634 702
rect 622 688 626 692
rect 654 758 658 762
rect 838 1058 842 1062
rect 822 998 826 1002
rect 814 978 818 982
rect 806 958 810 962
rect 950 1108 954 1112
rect 942 1098 946 1102
rect 970 1103 974 1107
rect 977 1103 981 1107
rect 918 1088 922 1092
rect 950 1088 954 1092
rect 1070 1448 1074 1452
rect 1102 1508 1106 1512
rect 1134 1488 1138 1492
rect 1102 1468 1106 1472
rect 1222 1538 1226 1542
rect 1190 1528 1194 1532
rect 1302 1538 1306 1542
rect 1294 1528 1298 1532
rect 1198 1518 1202 1522
rect 1254 1518 1258 1522
rect 1270 1508 1274 1512
rect 1174 1478 1178 1482
rect 1214 1478 1218 1482
rect 1238 1478 1242 1482
rect 1262 1478 1266 1482
rect 1246 1468 1250 1472
rect 1190 1459 1194 1463
rect 1198 1428 1202 1432
rect 1134 1358 1138 1362
rect 1254 1358 1258 1362
rect 1278 1428 1282 1432
rect 1278 1418 1282 1422
rect 1598 1668 1602 1672
rect 1446 1658 1450 1662
rect 1510 1658 1514 1662
rect 1526 1648 1530 1652
rect 1482 1603 1486 1607
rect 1489 1603 1493 1607
rect 1478 1588 1482 1592
rect 1446 1578 1450 1582
rect 1462 1558 1466 1562
rect 1550 1618 1554 1622
rect 1670 1658 1674 1662
rect 1646 1648 1650 1652
rect 1630 1638 1634 1642
rect 1614 1588 1618 1592
rect 1510 1558 1514 1562
rect 1342 1548 1346 1552
rect 1390 1548 1394 1552
rect 1398 1548 1402 1552
rect 1542 1548 1546 1552
rect 1326 1528 1330 1532
rect 1342 1528 1346 1532
rect 1382 1528 1386 1532
rect 1326 1518 1330 1522
rect 1350 1508 1354 1512
rect 1342 1468 1346 1472
rect 1446 1538 1450 1542
rect 1454 1488 1458 1492
rect 1470 1488 1474 1492
rect 1526 1538 1530 1542
rect 1518 1528 1522 1532
rect 1542 1528 1546 1532
rect 1566 1528 1570 1532
rect 1486 1478 1490 1482
rect 1358 1448 1362 1452
rect 1486 1458 1490 1462
rect 1662 1558 1666 1562
rect 1662 1538 1666 1542
rect 1630 1478 1634 1482
rect 1670 1478 1674 1482
rect 1614 1468 1618 1472
rect 1686 1698 1690 1702
rect 1702 1698 1706 1702
rect 1694 1648 1698 1652
rect 1718 1528 1722 1532
rect 1758 1578 1762 1582
rect 1790 1658 1794 1662
rect 1766 1558 1770 1562
rect 1758 1548 1762 1552
rect 1814 1548 1818 1552
rect 1718 1488 1722 1492
rect 1742 1538 1746 1542
rect 1774 1538 1778 1542
rect 1806 1538 1810 1542
rect 1926 1638 1930 1642
rect 1910 1578 1914 1582
rect 1854 1558 1858 1562
rect 1750 1488 1754 1492
rect 1822 1488 1826 1492
rect 1622 1458 1626 1462
rect 1734 1458 1738 1462
rect 1518 1448 1522 1452
rect 1630 1448 1634 1452
rect 1318 1438 1322 1442
rect 1422 1438 1426 1442
rect 1662 1448 1666 1452
rect 1702 1448 1706 1452
rect 1750 1448 1754 1452
rect 1710 1438 1714 1442
rect 1638 1428 1642 1432
rect 1318 1418 1322 1422
rect 1482 1403 1486 1407
rect 1489 1403 1493 1407
rect 1614 1388 1618 1392
rect 1310 1378 1314 1382
rect 1614 1378 1618 1382
rect 1374 1368 1378 1372
rect 1454 1368 1458 1372
rect 1494 1368 1498 1372
rect 1318 1358 1322 1362
rect 1342 1358 1346 1362
rect 1542 1358 1546 1362
rect 1574 1358 1578 1362
rect 1606 1358 1610 1362
rect 1054 1348 1058 1352
rect 1238 1348 1242 1352
rect 1334 1348 1338 1352
rect 1006 1248 1010 1252
rect 1030 1168 1034 1172
rect 1014 1118 1018 1122
rect 1102 1338 1106 1342
rect 1102 1308 1106 1312
rect 1110 1288 1114 1292
rect 1094 1268 1098 1272
rect 1206 1318 1210 1322
rect 1174 1288 1178 1292
rect 1198 1288 1202 1292
rect 1230 1268 1234 1272
rect 1270 1338 1274 1342
rect 1126 1258 1130 1262
rect 1262 1258 1266 1262
rect 1118 1238 1122 1242
rect 1102 1178 1106 1182
rect 1070 1148 1074 1152
rect 1094 1148 1098 1152
rect 1078 1138 1082 1142
rect 1030 1088 1034 1092
rect 1022 1078 1026 1082
rect 894 1059 898 1062
rect 894 1058 898 1059
rect 870 978 874 982
rect 990 1058 994 1062
rect 1046 1038 1050 1042
rect 1070 1038 1074 1042
rect 1030 1018 1034 1022
rect 990 998 994 1002
rect 742 948 746 952
rect 846 948 850 952
rect 718 818 722 822
rect 806 928 810 932
rect 814 918 818 922
rect 870 938 874 942
rect 1030 988 1034 992
rect 934 938 938 942
rect 878 928 882 932
rect 910 928 914 932
rect 790 858 794 862
rect 782 768 786 772
rect 774 758 778 762
rect 646 718 650 722
rect 702 718 706 722
rect 638 678 642 682
rect 598 658 602 662
rect 534 648 538 652
rect 590 648 594 652
rect 458 603 462 607
rect 465 603 469 607
rect 446 558 450 562
rect 454 558 458 562
rect 278 528 282 532
rect 302 528 306 532
rect 422 528 426 532
rect 278 498 282 502
rect 286 488 290 492
rect 302 488 306 492
rect 94 398 98 402
rect 94 388 98 392
rect 222 398 226 402
rect 142 348 146 352
rect 302 478 306 482
rect 334 498 338 502
rect 382 498 386 502
rect 406 498 410 502
rect 430 498 434 502
rect 390 488 394 492
rect 430 488 434 492
rect 510 578 514 582
rect 494 558 498 562
rect 518 558 522 562
rect 486 548 490 552
rect 510 548 514 552
rect 478 528 482 532
rect 486 488 490 492
rect 326 468 330 472
rect 374 468 378 472
rect 358 428 362 432
rect 286 358 290 362
rect 458 403 462 407
rect 465 403 469 407
rect 406 388 410 392
rect 390 358 394 362
rect 478 358 482 362
rect 502 358 506 362
rect 406 348 410 352
rect 454 348 458 352
rect 246 338 250 342
rect 326 338 330 342
rect 358 338 362 342
rect 422 338 426 342
rect 62 298 66 302
rect 110 298 114 302
rect 6 248 10 252
rect 38 248 42 252
rect 70 248 74 252
rect 78 238 82 242
rect 142 268 146 272
rect 126 258 130 262
rect 302 318 306 322
rect 350 288 354 292
rect 286 278 290 282
rect 206 248 210 252
rect 182 218 186 222
rect 110 158 114 162
rect 6 148 10 152
rect 86 148 90 152
rect 6 118 10 122
rect 38 118 42 122
rect 70 108 74 112
rect 174 138 178 142
rect 142 118 146 122
rect 134 108 138 112
rect 126 98 130 102
rect 126 88 130 92
rect 134 78 138 82
rect 166 78 170 82
rect 254 228 258 232
rect 302 228 306 232
rect 262 218 266 222
rect 382 308 386 312
rect 366 278 370 282
rect 406 278 410 282
rect 574 547 578 551
rect 582 538 586 542
rect 574 528 578 532
rect 558 478 562 482
rect 534 459 538 463
rect 526 388 530 392
rect 582 468 586 472
rect 518 348 522 352
rect 614 558 618 562
rect 670 698 674 702
rect 710 678 714 682
rect 694 668 698 672
rect 766 748 770 752
rect 766 738 770 742
rect 814 758 818 762
rect 814 748 818 752
rect 806 738 810 742
rect 734 728 738 732
rect 798 728 802 732
rect 782 718 786 722
rect 774 698 778 702
rect 790 688 794 692
rect 734 668 738 672
rect 766 668 770 672
rect 694 588 698 592
rect 670 547 674 551
rect 646 538 650 542
rect 686 488 690 492
rect 734 588 738 592
rect 726 568 730 572
rect 758 568 762 572
rect 766 558 770 562
rect 970 903 974 907
rect 977 903 981 907
rect 950 878 954 882
rect 862 828 866 832
rect 862 798 866 802
rect 830 778 834 782
rect 862 778 866 782
rect 1006 818 1010 822
rect 982 808 986 812
rect 838 758 842 762
rect 886 758 890 762
rect 918 758 922 762
rect 830 718 834 722
rect 990 798 994 802
rect 1102 1128 1106 1132
rect 1102 1118 1106 1122
rect 1102 1048 1106 1052
rect 1222 1248 1226 1252
rect 1318 1328 1322 1332
rect 1318 1298 1322 1302
rect 1366 1348 1370 1352
rect 1382 1348 1386 1352
rect 1414 1348 1418 1352
rect 1430 1348 1434 1352
rect 1454 1338 1458 1342
rect 1374 1328 1378 1332
rect 1438 1328 1442 1332
rect 1406 1318 1410 1322
rect 1454 1318 1458 1322
rect 1374 1308 1378 1312
rect 1398 1308 1402 1312
rect 1374 1268 1378 1272
rect 1518 1338 1522 1342
rect 1518 1328 1522 1332
rect 1478 1318 1482 1322
rect 1462 1308 1466 1312
rect 1470 1298 1474 1302
rect 1550 1338 1554 1342
rect 1574 1338 1578 1342
rect 1606 1338 1610 1342
rect 1606 1328 1610 1332
rect 1622 1328 1626 1332
rect 1534 1318 1538 1322
rect 1566 1318 1570 1322
rect 1502 1278 1506 1282
rect 1430 1268 1434 1272
rect 1294 1248 1298 1252
rect 1326 1238 1330 1242
rect 1278 1228 1282 1232
rect 1158 1218 1162 1222
rect 1262 1218 1266 1222
rect 1134 1168 1138 1172
rect 1126 1158 1130 1162
rect 1142 1148 1146 1152
rect 1134 1128 1138 1132
rect 1126 1108 1130 1112
rect 1238 1178 1242 1182
rect 1206 1138 1210 1142
rect 1254 1158 1258 1162
rect 1278 1178 1282 1182
rect 1310 1178 1314 1182
rect 1278 1168 1282 1172
rect 1246 1138 1250 1142
rect 1238 1118 1242 1122
rect 1230 1108 1234 1112
rect 1214 1098 1218 1102
rect 1166 1068 1170 1072
rect 1134 1058 1138 1062
rect 1118 988 1122 992
rect 1182 988 1186 992
rect 1118 978 1122 982
rect 1158 978 1162 982
rect 1078 938 1082 942
rect 1054 928 1058 932
rect 1070 888 1074 892
rect 1062 878 1066 882
rect 1046 868 1050 872
rect 1046 848 1050 852
rect 998 788 1002 792
rect 854 748 858 752
rect 878 748 882 752
rect 926 748 930 752
rect 982 748 986 752
rect 862 738 866 742
rect 862 708 866 712
rect 886 738 890 742
rect 966 718 970 722
rect 970 703 974 707
rect 977 703 981 707
rect 958 698 962 702
rect 1102 938 1106 942
rect 1134 938 1138 942
rect 1198 978 1202 982
rect 1174 938 1178 942
rect 1198 938 1202 942
rect 1150 918 1154 922
rect 1198 918 1202 922
rect 1134 888 1138 892
rect 1142 888 1146 892
rect 1110 868 1114 872
rect 1086 858 1090 862
rect 1078 808 1082 812
rect 1030 758 1034 762
rect 878 688 882 692
rect 886 688 890 692
rect 942 688 946 692
rect 974 688 978 692
rect 822 678 826 682
rect 878 678 882 682
rect 830 659 834 663
rect 934 678 938 682
rect 918 668 922 672
rect 942 668 946 672
rect 1038 668 1042 672
rect 878 658 882 662
rect 1174 878 1178 882
rect 1190 868 1194 872
rect 1262 1108 1266 1112
rect 1246 1088 1250 1092
rect 1222 1048 1226 1052
rect 1222 998 1226 1002
rect 1214 948 1218 952
rect 1214 878 1218 882
rect 1310 1168 1314 1172
rect 1366 1258 1370 1262
rect 1382 1248 1386 1252
rect 1390 1248 1394 1252
rect 1438 1258 1442 1262
rect 1462 1258 1466 1262
rect 1406 1208 1410 1212
rect 1358 1158 1362 1162
rect 1294 1148 1298 1152
rect 1310 1148 1314 1152
rect 1374 1148 1378 1152
rect 1294 1138 1298 1142
rect 1350 1138 1354 1142
rect 1302 1058 1306 1062
rect 1398 1138 1402 1142
rect 1374 1098 1378 1102
rect 1334 1088 1338 1092
rect 1358 1088 1362 1092
rect 1382 1078 1386 1082
rect 1350 1068 1354 1072
rect 1318 968 1322 972
rect 1334 968 1338 972
rect 1254 948 1258 952
rect 1310 938 1314 942
rect 1254 928 1258 932
rect 1278 918 1282 922
rect 1310 918 1314 922
rect 1318 918 1322 922
rect 1334 918 1338 922
rect 1238 888 1242 892
rect 1270 878 1274 882
rect 1430 1208 1434 1212
rect 1422 1148 1426 1152
rect 1478 1248 1482 1252
rect 1454 1208 1458 1212
rect 1482 1203 1486 1207
rect 1489 1203 1493 1207
rect 1502 1168 1506 1172
rect 1526 1268 1530 1272
rect 1550 1258 1554 1262
rect 1590 1278 1594 1282
rect 1574 1268 1578 1272
rect 1590 1248 1594 1252
rect 1558 1238 1562 1242
rect 1558 1158 1562 1162
rect 1566 1158 1570 1162
rect 1518 1148 1522 1152
rect 1494 1138 1498 1142
rect 1422 1088 1426 1092
rect 1414 1058 1418 1062
rect 1462 1098 1466 1102
rect 1470 1098 1474 1102
rect 1454 1088 1458 1092
rect 1542 1128 1546 1132
rect 1526 1118 1530 1122
rect 1526 1068 1530 1072
rect 1494 1058 1498 1062
rect 1550 1088 1554 1092
rect 1590 1098 1594 1102
rect 1566 1058 1570 1062
rect 1582 1058 1586 1062
rect 1510 1018 1514 1022
rect 1542 1018 1546 1022
rect 1482 1003 1486 1007
rect 1489 1003 1493 1007
rect 1430 988 1434 992
rect 1494 958 1498 962
rect 1534 988 1538 992
rect 1590 968 1594 972
rect 1622 1258 1626 1262
rect 1630 1258 1634 1262
rect 1806 1428 1810 1432
rect 1846 1448 1850 1452
rect 1902 1428 1906 1432
rect 1910 1378 1914 1382
rect 1646 1348 1650 1352
rect 1662 1348 1666 1352
rect 1686 1348 1690 1352
rect 1726 1351 1730 1352
rect 1726 1348 1730 1351
rect 1846 1348 1850 1352
rect 1654 1338 1658 1342
rect 1678 1338 1682 1342
rect 1726 1338 1730 1342
rect 1646 1328 1650 1332
rect 1670 1318 1674 1322
rect 1670 1278 1674 1282
rect 1606 1248 1610 1252
rect 1806 1338 1810 1342
rect 1830 1338 1834 1342
rect 1774 1258 1778 1262
rect 1718 1248 1722 1252
rect 1718 1238 1722 1242
rect 1654 1218 1658 1222
rect 1638 1188 1642 1192
rect 1686 1158 1690 1162
rect 1646 1147 1650 1151
rect 1670 1128 1674 1132
rect 1694 1128 1698 1132
rect 1646 1118 1650 1122
rect 1622 1098 1626 1102
rect 1606 1078 1610 1082
rect 1630 1078 1634 1082
rect 1670 1078 1674 1082
rect 1622 1068 1626 1072
rect 1646 1068 1650 1072
rect 1678 1068 1682 1072
rect 1686 1068 1690 1072
rect 1606 1058 1610 1062
rect 1630 1058 1634 1062
rect 1654 1058 1658 1062
rect 1598 948 1602 952
rect 1430 938 1434 942
rect 1662 938 1666 942
rect 1398 918 1402 922
rect 1430 908 1434 912
rect 1374 878 1378 882
rect 1422 878 1426 882
rect 1238 868 1242 872
rect 1326 868 1330 872
rect 1214 858 1218 862
rect 1262 858 1266 862
rect 1198 818 1202 822
rect 1142 788 1146 792
rect 1174 788 1178 792
rect 1214 788 1218 792
rect 1214 758 1218 762
rect 1270 758 1274 762
rect 1262 748 1266 752
rect 1110 738 1114 742
rect 1166 738 1170 742
rect 1094 728 1098 732
rect 1086 718 1090 722
rect 1110 718 1114 722
rect 1070 668 1074 672
rect 1166 688 1170 692
rect 1134 678 1138 682
rect 1238 738 1242 742
rect 1286 738 1290 742
rect 1254 728 1258 732
rect 1278 728 1282 732
rect 1222 638 1226 642
rect 1374 868 1378 872
rect 1454 878 1458 882
rect 1726 1158 1730 1162
rect 1734 1148 1738 1152
rect 1718 1108 1722 1112
rect 1790 1248 1794 1252
rect 1790 1218 1794 1222
rect 1750 1168 1754 1172
rect 1774 1168 1778 1172
rect 1798 1148 1802 1152
rect 1742 1138 1746 1142
rect 1886 1288 1890 1292
rect 1838 1278 1842 1282
rect 1918 1268 1922 1272
rect 1886 1258 1890 1262
rect 1918 1258 1922 1262
rect 1830 1238 1834 1242
rect 1894 1238 1898 1242
rect 1822 1178 1826 1182
rect 1862 1178 1866 1182
rect 1838 1158 1842 1162
rect 1862 1158 1866 1162
rect 1830 1148 1834 1152
rect 1854 1148 1858 1152
rect 1766 1128 1770 1132
rect 1806 1128 1810 1132
rect 1854 1128 1858 1132
rect 1878 1158 1882 1162
rect 1926 1248 1930 1252
rect 1934 1238 1938 1242
rect 1894 1148 1898 1152
rect 1886 1138 1890 1142
rect 1902 1128 1906 1132
rect 1950 1548 1954 1552
rect 1950 1348 1954 1352
rect 1950 1268 1954 1272
rect 1918 1088 1922 1092
rect 1942 1088 1946 1092
rect 1902 1068 1906 1072
rect 1822 1058 1826 1062
rect 1750 1048 1754 1052
rect 1806 988 1810 992
rect 1838 988 1842 992
rect 1766 958 1770 962
rect 1742 948 1746 952
rect 1790 948 1794 952
rect 1694 938 1698 942
rect 1726 938 1730 942
rect 1678 908 1682 912
rect 1502 868 1506 872
rect 1534 868 1538 872
rect 1390 858 1394 862
rect 1406 858 1410 862
rect 1382 848 1386 852
rect 1374 838 1378 842
rect 1482 803 1486 807
rect 1489 803 1493 807
rect 1598 898 1602 902
rect 1718 918 1722 922
rect 1726 918 1730 922
rect 1862 947 1866 951
rect 1942 948 1946 952
rect 1910 918 1914 922
rect 1918 908 1922 912
rect 1838 888 1842 892
rect 1742 878 1746 882
rect 1758 878 1762 882
rect 1814 878 1818 882
rect 1638 868 1642 872
rect 1694 868 1698 872
rect 1574 858 1578 862
rect 1590 858 1594 862
rect 1606 858 1610 862
rect 1622 818 1626 822
rect 1654 858 1658 862
rect 1662 848 1666 852
rect 1678 848 1682 852
rect 1646 828 1650 832
rect 1654 818 1658 822
rect 1374 778 1378 782
rect 1686 838 1690 842
rect 1710 838 1714 842
rect 1750 848 1754 852
rect 1734 828 1738 832
rect 1782 828 1786 832
rect 1662 768 1666 772
rect 1646 758 1650 762
rect 1662 758 1666 762
rect 1590 748 1594 752
rect 1646 748 1650 752
rect 1342 738 1346 742
rect 1366 738 1370 742
rect 1374 738 1378 742
rect 1398 698 1402 702
rect 1334 688 1338 692
rect 1350 658 1354 662
rect 1246 638 1250 642
rect 1462 738 1466 742
rect 1478 698 1482 702
rect 1422 658 1426 662
rect 1470 658 1474 662
rect 1238 628 1242 632
rect 1406 628 1410 632
rect 1054 568 1058 572
rect 1102 568 1106 572
rect 1158 568 1162 572
rect 806 558 810 562
rect 838 558 842 562
rect 862 558 866 562
rect 870 558 874 562
rect 1038 558 1042 562
rect 1054 558 1058 562
rect 710 548 714 552
rect 758 548 762 552
rect 878 548 882 552
rect 1086 548 1090 552
rect 726 538 730 542
rect 774 538 778 542
rect 838 538 842 542
rect 878 538 882 542
rect 726 528 730 532
rect 838 528 842 532
rect 862 528 866 532
rect 870 528 874 532
rect 902 528 906 532
rect 934 528 938 532
rect 710 518 714 522
rect 638 478 642 482
rect 686 478 690 482
rect 790 488 794 492
rect 806 478 810 482
rect 830 478 834 482
rect 822 468 826 472
rect 742 458 746 462
rect 694 358 698 362
rect 678 348 682 352
rect 494 338 498 342
rect 510 338 514 342
rect 502 328 506 332
rect 534 328 538 332
rect 430 308 434 312
rect 478 288 482 292
rect 846 438 850 442
rect 886 498 890 502
rect 902 478 906 482
rect 918 468 922 472
rect 902 458 906 462
rect 926 458 930 462
rect 950 458 954 462
rect 910 448 914 452
rect 886 388 890 392
rect 918 358 922 362
rect 854 348 858 352
rect 726 338 730 342
rect 750 338 754 342
rect 678 328 682 332
rect 654 318 658 322
rect 382 258 386 262
rect 510 238 514 242
rect 406 228 410 232
rect 206 168 210 172
rect 238 168 242 172
rect 458 203 462 207
rect 465 203 469 207
rect 470 168 474 172
rect 486 168 490 172
rect 414 158 418 162
rect 190 148 194 152
rect 238 148 242 152
rect 294 148 298 152
rect 318 148 322 152
rect 350 148 354 152
rect 262 138 266 142
rect 286 138 290 142
rect 230 118 234 122
rect 270 118 274 122
rect 302 118 306 122
rect 302 108 306 112
rect 270 98 274 102
rect 214 88 218 92
rect 206 78 210 82
rect 110 68 114 72
rect 158 68 162 72
rect 174 68 178 72
rect 310 88 314 92
rect 238 78 242 82
rect 294 78 298 82
rect 326 78 330 82
rect 230 68 234 72
rect 38 58 42 62
rect 150 58 154 62
rect 166 58 170 62
rect 54 48 58 52
rect 142 48 146 52
rect 158 48 162 52
rect 198 48 202 52
rect 598 158 602 162
rect 558 148 562 152
rect 430 128 434 132
rect 454 108 458 112
rect 462 108 466 112
rect 414 98 418 102
rect 358 88 362 92
rect 342 68 346 72
rect 502 118 506 122
rect 550 118 554 122
rect 470 88 474 92
rect 486 78 490 82
rect 518 68 522 72
rect 414 48 418 52
rect 494 48 498 52
rect 510 48 514 52
rect 598 138 602 142
rect 574 128 578 132
rect 614 128 618 132
rect 606 88 610 92
rect 686 288 690 292
rect 790 328 794 332
rect 766 278 770 282
rect 750 258 754 262
rect 774 258 778 262
rect 694 248 698 252
rect 1030 528 1034 532
rect 982 518 986 522
rect 970 503 974 507
rect 977 503 981 507
rect 1006 488 1010 492
rect 990 448 994 452
rect 1086 538 1090 542
rect 1094 538 1098 542
rect 1062 478 1066 482
rect 1046 468 1050 472
rect 1070 468 1074 472
rect 1014 458 1018 462
rect 958 388 962 392
rect 974 388 978 392
rect 990 338 994 342
rect 1014 340 1018 344
rect 1118 558 1122 562
rect 1126 548 1130 552
rect 1142 548 1146 552
rect 1174 548 1178 552
rect 1214 548 1218 552
rect 1630 738 1634 742
rect 1550 728 1554 732
rect 1526 718 1530 722
rect 1734 768 1738 772
rect 1686 758 1690 762
rect 1702 758 1706 762
rect 1646 738 1650 742
rect 1670 738 1674 742
rect 1638 708 1642 712
rect 1550 688 1554 692
rect 1606 678 1610 682
rect 1694 728 1698 732
rect 1654 718 1658 722
rect 1678 718 1682 722
rect 1662 688 1666 692
rect 1694 678 1698 682
rect 1550 668 1554 672
rect 1590 668 1594 672
rect 1630 668 1634 672
rect 1646 668 1650 672
rect 1662 668 1666 672
rect 1542 658 1546 662
rect 1646 648 1650 652
rect 1598 638 1602 642
rect 1482 603 1486 607
rect 1489 603 1493 607
rect 1398 578 1402 582
rect 1406 578 1410 582
rect 1494 578 1498 582
rect 1182 538 1186 542
rect 1198 538 1202 542
rect 1206 538 1210 542
rect 1302 538 1306 542
rect 1134 528 1138 532
rect 1150 528 1154 532
rect 1118 508 1122 512
rect 1142 518 1146 522
rect 1102 438 1106 442
rect 1062 388 1066 392
rect 1118 368 1122 372
rect 1038 338 1042 342
rect 1054 338 1058 342
rect 950 328 954 332
rect 970 303 974 307
rect 977 303 981 307
rect 958 278 962 282
rect 1038 328 1042 332
rect 1190 488 1194 492
rect 1198 468 1202 472
rect 1150 458 1154 462
rect 1158 448 1162 452
rect 1182 368 1186 372
rect 1134 338 1138 342
rect 1126 328 1130 332
rect 1086 308 1090 312
rect 1054 268 1058 272
rect 734 238 738 242
rect 758 238 762 242
rect 782 238 786 242
rect 814 238 818 242
rect 718 228 722 232
rect 742 228 746 232
rect 790 218 794 222
rect 806 218 810 222
rect 758 178 762 182
rect 694 168 698 172
rect 670 158 674 162
rect 750 158 754 162
rect 774 158 778 162
rect 646 138 650 142
rect 638 108 642 112
rect 622 98 626 102
rect 590 68 594 72
rect 614 68 618 72
rect 598 58 602 62
rect 638 58 642 62
rect 550 48 554 52
rect 254 38 258 42
rect 294 38 298 42
rect 534 38 538 42
rect 458 3 462 7
rect 465 3 469 7
rect 670 98 674 102
rect 870 218 874 222
rect 918 218 922 222
rect 1022 208 1026 212
rect 1086 198 1090 202
rect 846 188 850 192
rect 934 188 938 192
rect 878 178 882 182
rect 814 158 818 162
rect 886 148 890 152
rect 814 138 818 142
rect 838 138 842 142
rect 870 138 874 142
rect 782 128 786 132
rect 750 88 754 92
rect 822 128 826 132
rect 790 118 794 122
rect 814 118 818 122
rect 822 118 826 122
rect 798 108 802 112
rect 822 108 826 112
rect 814 98 818 102
rect 790 88 794 92
rect 862 98 866 102
rect 918 138 922 142
rect 926 128 930 132
rect 1006 138 1010 142
rect 902 118 906 122
rect 990 118 994 122
rect 1006 118 1010 122
rect 970 103 974 107
rect 977 103 981 107
rect 862 88 866 92
rect 918 88 922 92
rect 798 78 802 82
rect 926 78 930 82
rect 774 68 778 72
rect 790 68 794 72
rect 854 68 858 72
rect 878 68 882 72
rect 1046 118 1050 122
rect 1190 358 1194 362
rect 1238 518 1242 522
rect 1366 528 1370 532
rect 1478 568 1482 572
rect 1390 508 1394 512
rect 1374 488 1378 492
rect 1398 488 1402 492
rect 1454 548 1458 552
rect 1470 548 1474 552
rect 1526 548 1530 552
rect 1590 538 1594 542
rect 1518 528 1522 532
rect 1438 478 1442 482
rect 1246 468 1250 472
rect 1262 468 1266 472
rect 1302 468 1306 472
rect 1350 468 1354 472
rect 1454 468 1458 472
rect 1510 468 1514 472
rect 1214 368 1218 372
rect 1238 358 1242 362
rect 1334 458 1338 462
rect 1558 528 1562 532
rect 1566 518 1570 522
rect 1526 488 1530 492
rect 1534 478 1538 482
rect 1630 638 1634 642
rect 1606 628 1610 632
rect 1622 628 1626 632
rect 1638 578 1642 582
rect 1630 558 1634 562
rect 1606 548 1610 552
rect 1614 528 1618 532
rect 1598 508 1602 512
rect 1590 488 1594 492
rect 1526 458 1530 462
rect 1550 458 1554 462
rect 1558 458 1562 462
rect 1574 458 1578 462
rect 1582 458 1586 462
rect 1566 438 1570 442
rect 1550 428 1554 432
rect 1482 403 1486 407
rect 1489 403 1493 407
rect 1206 348 1210 352
rect 1390 348 1394 352
rect 1518 348 1522 352
rect 1446 338 1450 342
rect 1206 308 1210 312
rect 1238 308 1242 312
rect 1294 308 1298 312
rect 1350 308 1354 312
rect 1286 268 1290 272
rect 1390 268 1394 272
rect 1494 258 1498 262
rect 1118 208 1122 212
rect 1110 198 1114 202
rect 1094 148 1098 152
rect 1102 148 1106 152
rect 1078 138 1082 142
rect 1038 108 1042 112
rect 1054 108 1058 112
rect 1062 108 1066 112
rect 1006 88 1010 92
rect 1038 88 1042 92
rect 1334 248 1338 252
rect 1374 238 1378 242
rect 1454 238 1458 242
rect 1174 198 1178 202
rect 1278 158 1282 162
rect 1342 158 1346 162
rect 1398 158 1402 162
rect 1150 108 1154 112
rect 1158 98 1162 102
rect 1254 148 1258 152
rect 1190 138 1194 142
rect 1206 118 1210 122
rect 1206 98 1210 102
rect 1150 78 1154 82
rect 998 68 1002 72
rect 1006 68 1010 72
rect 1022 68 1026 72
rect 1070 68 1074 72
rect 1118 68 1122 72
rect 1134 68 1138 72
rect 982 58 986 62
rect 1046 58 1050 62
rect 1086 58 1090 62
rect 1214 88 1218 92
rect 1230 88 1234 92
rect 1230 78 1234 82
rect 1246 78 1250 82
rect 1198 58 1202 62
rect 854 48 858 52
rect 878 48 882 52
rect 1318 148 1322 152
rect 1310 138 1314 142
rect 1262 88 1266 92
rect 1294 78 1298 82
rect 1270 58 1274 62
rect 1278 58 1282 62
rect 1430 188 1434 192
rect 1366 148 1370 152
rect 1414 148 1418 152
rect 1438 148 1442 152
rect 1486 218 1490 222
rect 1482 203 1486 207
rect 1489 203 1493 207
rect 1622 498 1626 502
rect 1614 438 1618 442
rect 1574 428 1578 432
rect 1582 328 1586 332
rect 1550 288 1554 292
rect 1574 248 1578 252
rect 1518 188 1522 192
rect 1542 158 1546 162
rect 1358 118 1362 122
rect 1390 138 1394 142
rect 1422 138 1426 142
rect 1406 118 1410 122
rect 1398 108 1402 112
rect 1350 98 1354 102
rect 1374 98 1378 102
rect 1390 98 1394 102
rect 1366 88 1370 92
rect 1414 88 1418 92
rect 1550 148 1554 152
rect 1654 518 1658 522
rect 1646 488 1650 492
rect 1702 658 1706 662
rect 1694 638 1698 642
rect 1718 628 1722 632
rect 1670 578 1674 582
rect 1702 578 1706 582
rect 1694 558 1698 562
rect 1710 558 1714 562
rect 1718 558 1722 562
rect 1670 548 1674 552
rect 1782 768 1786 772
rect 1742 748 1746 752
rect 1758 728 1762 732
rect 1734 698 1738 702
rect 1774 708 1778 712
rect 1838 848 1842 852
rect 1806 768 1810 772
rect 1798 758 1802 762
rect 1950 908 1954 912
rect 1950 868 1954 872
rect 1862 828 1866 832
rect 1854 748 1858 752
rect 1790 688 1794 692
rect 1838 688 1842 692
rect 1806 678 1810 682
rect 1926 698 1930 702
rect 1878 688 1882 692
rect 1822 668 1826 672
rect 1870 668 1874 672
rect 1742 658 1746 662
rect 1750 658 1754 662
rect 1782 658 1786 662
rect 1734 648 1738 652
rect 1910 648 1914 652
rect 1782 568 1786 572
rect 1862 568 1866 572
rect 1798 558 1802 562
rect 1758 548 1762 552
rect 1774 548 1778 552
rect 1798 548 1802 552
rect 1678 538 1682 542
rect 1710 538 1714 542
rect 1726 538 1730 542
rect 1766 538 1770 542
rect 1790 538 1794 542
rect 1638 459 1642 463
rect 1726 528 1730 532
rect 1686 498 1690 502
rect 1718 498 1722 502
rect 1694 478 1698 482
rect 1686 468 1690 472
rect 1750 468 1754 472
rect 1710 458 1714 462
rect 1686 448 1690 452
rect 1662 438 1666 442
rect 1934 688 1938 692
rect 1950 668 1954 672
rect 1934 598 1938 602
rect 1822 538 1826 542
rect 1806 498 1810 502
rect 1806 488 1810 492
rect 1798 458 1802 462
rect 1782 428 1786 432
rect 1622 348 1626 352
rect 1686 348 1690 352
rect 1742 348 1746 352
rect 1750 348 1754 352
rect 1734 338 1738 342
rect 1678 298 1682 302
rect 1622 288 1626 292
rect 1654 288 1658 292
rect 1670 288 1674 292
rect 1702 298 1706 302
rect 1670 278 1674 282
rect 1686 278 1690 282
rect 1598 258 1602 262
rect 1550 138 1554 142
rect 1542 128 1546 132
rect 1446 88 1450 92
rect 1502 98 1506 102
rect 1454 78 1458 82
rect 1582 118 1586 122
rect 1622 118 1626 122
rect 1582 88 1586 92
rect 1622 88 1626 92
rect 1774 288 1778 292
rect 1790 288 1794 292
rect 1822 288 1826 292
rect 1718 258 1722 262
rect 1806 258 1810 262
rect 1734 188 1738 192
rect 1774 188 1778 192
rect 1766 158 1770 162
rect 1686 148 1690 152
rect 1726 148 1730 152
rect 1646 138 1650 142
rect 1694 138 1698 142
rect 1670 118 1674 122
rect 1670 88 1674 92
rect 1630 78 1634 82
rect 1590 68 1594 72
rect 1390 58 1394 62
rect 1574 58 1578 62
rect 1630 58 1634 62
rect 1678 58 1682 62
rect 1702 118 1706 122
rect 1934 528 1938 532
rect 1854 468 1858 472
rect 1846 458 1850 462
rect 1798 158 1802 162
rect 1782 138 1786 142
rect 1814 128 1818 132
rect 1726 118 1730 122
rect 1774 118 1778 122
rect 1806 118 1810 122
rect 1758 88 1762 92
rect 1838 148 1842 152
rect 1886 158 1890 162
rect 1878 151 1882 152
rect 1878 148 1882 151
rect 1838 138 1842 142
rect 1830 118 1834 122
rect 1718 78 1722 82
rect 1782 78 1786 82
rect 1854 78 1858 82
rect 1758 68 1762 72
rect 1942 128 1946 132
rect 1182 48 1186 52
rect 1222 48 1226 52
rect 1230 48 1234 52
rect 1262 48 1266 52
rect 1334 48 1338 52
rect 1822 48 1826 52
rect 846 38 850 42
rect 1030 38 1034 42
rect 1070 38 1074 42
rect 1630 38 1634 42
rect 766 18 770 22
rect 1482 3 1486 7
rect 1489 3 1493 7
<< metal3 >>
rect 968 1703 970 1707
rect 974 1703 977 1707
rect 982 1703 984 1707
rect 1066 1698 1070 1701
rect 1154 1698 1158 1701
rect 1322 1698 1326 1701
rect 1514 1698 1526 1701
rect 1690 1698 1702 1701
rect 1062 1688 1078 1691
rect 1062 1682 1065 1688
rect 98 1678 126 1681
rect 210 1678 214 1681
rect 410 1678 430 1681
rect 434 1678 622 1681
rect 1154 1678 1382 1681
rect 1386 1678 1446 1681
rect -26 1671 -22 1672
rect 6 1671 9 1678
rect -26 1668 9 1671
rect 62 1671 65 1678
rect 26 1668 65 1671
rect 134 1671 137 1678
rect 114 1668 129 1671
rect 134 1668 182 1671
rect 626 1668 694 1671
rect 1274 1668 1390 1671
rect 1394 1668 1454 1671
rect 1474 1668 1510 1671
rect 58 1658 86 1661
rect 126 1661 129 1668
rect 126 1658 166 1661
rect 430 1661 433 1668
rect 294 1658 433 1661
rect 438 1661 441 1668
rect 438 1658 478 1661
rect 574 1661 577 1668
rect 482 1658 489 1661
rect 574 1658 614 1661
rect 618 1658 662 1661
rect 874 1658 894 1661
rect 974 1661 977 1668
rect 974 1658 1006 1661
rect 1010 1658 1118 1661
rect 1154 1658 1158 1661
rect 1450 1658 1510 1661
rect 1598 1661 1601 1668
rect 1598 1658 1670 1661
rect 1694 1658 1790 1661
rect -26 1651 -22 1652
rect -26 1648 30 1651
rect 118 1651 121 1658
rect 294 1652 297 1658
rect 390 1652 393 1658
rect 1694 1652 1697 1658
rect 118 1648 150 1651
rect 498 1648 726 1651
rect 1042 1648 1118 1651
rect 1530 1648 1646 1651
rect 1022 1642 1025 1648
rect 74 1638 102 1641
rect 106 1638 142 1641
rect 146 1638 262 1641
rect 610 1638 646 1641
rect 1634 1638 1926 1641
rect 810 1628 822 1631
rect 826 1628 942 1631
rect 1322 1628 1326 1631
rect 1246 1622 1249 1628
rect 242 1618 254 1621
rect 258 1618 318 1621
rect 322 1618 470 1621
rect 522 1618 630 1621
rect 866 1618 918 1621
rect 922 1618 1078 1621
rect 1082 1618 1110 1621
rect 1554 1618 1654 1621
rect 1066 1608 1070 1611
rect 456 1603 458 1607
rect 462 1603 465 1607
rect 470 1603 472 1607
rect 1480 1603 1482 1607
rect 1486 1603 1489 1607
rect 1494 1603 1496 1607
rect 1194 1598 1270 1601
rect 1274 1598 1294 1601
rect 570 1588 1478 1591
rect 1482 1588 1614 1591
rect 442 1578 446 1581
rect 1218 1578 1310 1581
rect 1314 1578 1446 1581
rect 1762 1578 1910 1581
rect 994 1568 1030 1571
rect 378 1558 550 1561
rect 730 1558 910 1561
rect 954 1558 1014 1561
rect 1186 1558 1238 1561
rect 1666 1558 1766 1561
rect 170 1548 198 1551
rect 358 1551 361 1558
rect 358 1548 414 1551
rect 774 1548 870 1551
rect 962 1548 998 1551
rect 1026 1548 1086 1551
rect 1154 1548 1214 1551
rect 1266 1548 1278 1551
rect 1286 1551 1289 1558
rect 1286 1548 1305 1551
rect 1346 1548 1390 1551
rect 1394 1548 1398 1551
rect 1462 1551 1465 1558
rect 1510 1551 1513 1558
rect 1462 1548 1513 1551
rect 1746 1548 1758 1551
rect 1854 1551 1857 1558
rect 1818 1548 1857 1551
rect 1982 1551 1986 1552
rect 1954 1548 1986 1551
rect 774 1542 777 1548
rect 146 1538 190 1541
rect 194 1538 238 1541
rect 242 1538 286 1541
rect 290 1538 510 1541
rect 598 1538 606 1541
rect 850 1538 926 1541
rect 958 1541 961 1548
rect 930 1538 961 1541
rect 1262 1541 1265 1548
rect 1226 1538 1265 1541
rect 1302 1542 1305 1548
rect 1450 1538 1526 1541
rect 1542 1541 1545 1548
rect 1742 1542 1745 1548
rect 1530 1538 1662 1541
rect 1778 1538 1806 1541
rect 598 1532 601 1538
rect 698 1528 774 1531
rect 906 1528 958 1531
rect 962 1528 966 1531
rect 1018 1528 1038 1531
rect 1090 1528 1190 1531
rect 1298 1528 1326 1531
rect 1346 1528 1382 1531
rect 1522 1528 1542 1531
rect 1546 1528 1566 1531
rect 1658 1528 1718 1531
rect 306 1518 430 1521
rect 434 1518 470 1521
rect 530 1518 582 1521
rect 586 1518 606 1521
rect 1202 1518 1254 1521
rect 1330 1518 1353 1521
rect 1350 1512 1353 1518
rect 210 1508 566 1511
rect 578 1508 614 1511
rect 618 1508 670 1511
rect 714 1508 806 1511
rect 810 1508 814 1511
rect 1106 1508 1270 1511
rect 968 1503 970 1507
rect 974 1503 977 1507
rect 982 1503 984 1507
rect 314 1498 422 1501
rect 514 1498 686 1501
rect 914 1488 1046 1491
rect 1050 1488 1134 1491
rect 1138 1488 1454 1491
rect 1474 1488 1718 1491
rect 1722 1488 1750 1491
rect 1754 1488 1822 1491
rect 242 1478 334 1481
rect 534 1481 537 1488
rect 338 1478 537 1481
rect 710 1481 713 1488
rect 634 1478 713 1481
rect 826 1478 846 1481
rect 850 1478 1022 1481
rect 1026 1478 1030 1481
rect 1042 1478 1174 1481
rect 1234 1478 1238 1481
rect 1266 1478 1486 1481
rect 1626 1478 1630 1481
rect 370 1468 398 1471
rect 410 1468 422 1471
rect 442 1468 518 1471
rect 522 1468 670 1471
rect 786 1468 862 1471
rect 890 1468 993 1471
rect 62 1461 65 1468
rect 110 1461 113 1468
rect 62 1458 113 1461
rect 118 1461 121 1468
rect 118 1458 142 1461
rect 146 1458 153 1461
rect 258 1458 374 1461
rect 418 1458 446 1461
rect 514 1458 526 1461
rect 578 1458 590 1461
rect 990 1462 993 1468
rect 1214 1471 1217 1478
rect 1214 1468 1246 1471
rect 1250 1468 1342 1471
rect 1670 1471 1673 1478
rect 1618 1468 1673 1471
rect 802 1459 838 1461
rect 798 1458 838 1459
rect 874 1458 918 1461
rect 946 1458 966 1461
rect 1102 1461 1105 1468
rect 994 1458 1073 1461
rect 1102 1459 1190 1461
rect 1194 1459 1230 1461
rect 1102 1458 1230 1459
rect 1490 1458 1622 1461
rect 1626 1458 1734 1461
rect 1070 1452 1073 1458
rect 378 1448 558 1451
rect 562 1448 718 1451
rect 722 1448 886 1451
rect 946 1448 958 1451
rect 1074 1448 1246 1451
rect 1250 1448 1358 1451
rect 1362 1448 1518 1451
rect 1626 1448 1630 1451
rect 1654 1448 1662 1451
rect 1666 1448 1702 1451
rect 1710 1448 1750 1451
rect 1754 1448 1846 1451
rect 1710 1442 1713 1448
rect 18 1438 126 1441
rect 130 1438 134 1441
rect 394 1438 422 1441
rect 426 1438 518 1441
rect 634 1438 806 1441
rect 834 1438 854 1441
rect 1226 1438 1318 1441
rect 1322 1438 1422 1441
rect 386 1428 638 1431
rect 738 1428 862 1431
rect 906 1428 934 1431
rect 1202 1428 1278 1431
rect 1386 1428 1638 1431
rect 1642 1428 1806 1431
rect 1810 1428 1902 1431
rect 186 1418 270 1421
rect 754 1418 814 1421
rect 1282 1418 1318 1421
rect 666 1408 902 1411
rect 456 1403 458 1407
rect 462 1403 465 1407
rect 470 1403 472 1407
rect 1480 1403 1482 1407
rect 1486 1403 1489 1407
rect 1494 1403 1496 1407
rect 74 1398 254 1401
rect 258 1398 286 1401
rect 522 1398 542 1401
rect 546 1398 574 1401
rect 362 1388 446 1391
rect 450 1388 630 1391
rect 1594 1388 1614 1391
rect 706 1378 790 1381
rect 794 1378 1006 1381
rect 1122 1378 1310 1381
rect 1314 1378 1614 1381
rect 1618 1378 1734 1381
rect 162 1368 382 1371
rect 666 1368 710 1371
rect 738 1368 742 1371
rect 1318 1368 1374 1371
rect 1458 1368 1494 1371
rect 1910 1371 1913 1378
rect 1982 1371 1986 1372
rect 1910 1368 1986 1371
rect 10 1358 190 1361
rect 194 1358 230 1361
rect 274 1358 278 1361
rect 378 1358 438 1361
rect 570 1358 614 1361
rect 618 1358 638 1361
rect 718 1361 721 1368
rect 1318 1362 1321 1368
rect 642 1358 721 1361
rect 1138 1358 1254 1361
rect 1346 1358 1542 1361
rect 1546 1358 1574 1361
rect 1578 1358 1606 1361
rect 122 1348 126 1351
rect 130 1348 225 1351
rect 306 1348 318 1351
rect 634 1348 678 1351
rect 682 1348 694 1351
rect 714 1348 758 1351
rect 930 1348 934 1351
rect 1014 1351 1017 1358
rect 970 1348 1017 1351
rect 1058 1348 1230 1351
rect 1234 1348 1238 1351
rect 1270 1348 1302 1351
rect 1338 1348 1366 1351
rect 1370 1348 1382 1351
rect 1386 1348 1414 1351
rect 1650 1348 1654 1351
rect 1666 1348 1686 1351
rect 1730 1348 1846 1351
rect 1982 1351 1986 1352
rect 1954 1348 1986 1351
rect 222 1342 225 1348
rect 66 1338 134 1341
rect 138 1338 198 1341
rect 330 1338 350 1341
rect 426 1338 438 1341
rect 562 1338 566 1341
rect 594 1338 614 1341
rect 658 1338 726 1341
rect 846 1341 849 1348
rect 1270 1342 1273 1348
rect 738 1338 849 1341
rect 858 1338 918 1341
rect 922 1338 1102 1341
rect 1374 1338 1414 1341
rect 1430 1341 1433 1348
rect 1430 1338 1454 1341
rect 1522 1338 1550 1341
rect 1578 1338 1582 1341
rect 1610 1338 1654 1341
rect 1682 1338 1726 1341
rect 1810 1338 1830 1341
rect 1374 1332 1377 1338
rect 146 1328 190 1331
rect 194 1328 206 1331
rect 218 1328 246 1331
rect 378 1328 390 1331
rect 714 1328 750 1331
rect 762 1328 1318 1331
rect 1442 1328 1518 1331
rect 1610 1328 1622 1331
rect 1650 1328 1673 1331
rect 302 1321 305 1328
rect 1670 1322 1673 1328
rect 242 1318 305 1321
rect 530 1318 542 1321
rect 546 1318 654 1321
rect 690 1318 718 1321
rect 842 1318 1206 1321
rect 1410 1318 1454 1321
rect 1482 1318 1534 1321
rect 1538 1318 1566 1321
rect 290 1308 342 1311
rect 378 1308 430 1311
rect 570 1308 638 1311
rect 642 1308 878 1311
rect 890 1308 894 1311
rect 1106 1308 1374 1311
rect 1402 1308 1462 1311
rect 968 1303 970 1307
rect 974 1303 977 1307
rect 982 1303 984 1307
rect 66 1298 406 1301
rect 514 1298 574 1301
rect 842 1298 846 1301
rect 1322 1298 1470 1301
rect 302 1288 430 1291
rect 434 1288 478 1291
rect 482 1288 486 1291
rect 730 1288 830 1291
rect 1114 1288 1174 1291
rect 302 1282 305 1288
rect 346 1278 422 1281
rect 518 1281 521 1288
rect 426 1278 441 1281
rect 518 1278 598 1281
rect 810 1278 838 1281
rect 1174 1281 1177 1288
rect 1198 1281 1201 1288
rect 1174 1278 1201 1281
rect 1506 1278 1590 1281
rect 1886 1281 1889 1288
rect 1842 1278 1889 1281
rect 86 1271 89 1278
rect 438 1272 441 1278
rect 86 1268 142 1271
rect 274 1268 294 1271
rect 298 1268 302 1271
rect 338 1268 382 1271
rect 718 1271 721 1278
rect 530 1268 721 1271
rect 1098 1268 1222 1271
rect 1226 1268 1230 1271
rect 1378 1268 1430 1271
rect 1578 1268 1598 1271
rect 1670 1271 1673 1278
rect 1602 1268 1673 1271
rect 1922 1268 1934 1271
rect 1938 1268 1950 1271
rect 154 1258 158 1261
rect 166 1261 169 1268
rect 166 1258 238 1261
rect 338 1258 526 1261
rect 562 1258 598 1261
rect 674 1258 694 1261
rect 798 1261 801 1268
rect 798 1258 854 1261
rect 874 1258 958 1261
rect 1130 1258 1262 1261
rect 1370 1258 1438 1261
rect 1526 1261 1529 1268
rect 1466 1258 1529 1261
rect 1554 1258 1622 1261
rect 1634 1258 1774 1261
rect 1890 1258 1918 1261
rect 378 1248 382 1251
rect 402 1248 406 1251
rect 426 1248 502 1251
rect 630 1251 633 1258
rect 630 1248 678 1251
rect 682 1248 726 1251
rect 738 1248 801 1251
rect 834 1248 886 1251
rect 1010 1248 1222 1251
rect 1226 1248 1294 1251
rect 1394 1248 1398 1251
rect 1482 1248 1561 1251
rect 1594 1248 1606 1251
rect 1610 1248 1718 1251
rect 1722 1248 1790 1251
rect 1982 1251 1986 1252
rect 1930 1248 1986 1251
rect 18 1238 86 1241
rect 90 1238 334 1241
rect 394 1238 406 1241
rect 558 1241 561 1248
rect 798 1242 801 1248
rect 1382 1242 1385 1248
rect 1558 1242 1561 1248
rect 558 1238 590 1241
rect 602 1238 782 1241
rect 1122 1238 1326 1241
rect 1658 1238 1718 1241
rect 1722 1238 1830 1241
rect 1898 1238 1934 1241
rect 578 1228 670 1231
rect 698 1228 766 1231
rect 910 1231 913 1238
rect 770 1228 913 1231
rect 1282 1228 1286 1231
rect 1162 1218 1262 1221
rect 1266 1218 1654 1221
rect 1658 1218 1742 1221
rect 1746 1218 1790 1221
rect 482 1208 550 1211
rect 1410 1208 1430 1211
rect 1434 1208 1454 1211
rect 456 1203 458 1207
rect 462 1203 465 1207
rect 470 1203 472 1207
rect 1480 1203 1482 1207
rect 1486 1203 1489 1207
rect 1494 1203 1496 1207
rect 482 1198 566 1201
rect 818 1198 822 1201
rect 1402 1188 1638 1191
rect 518 1181 521 1188
rect 402 1178 521 1181
rect 762 1178 870 1181
rect 1106 1178 1238 1181
rect 1242 1178 1278 1181
rect 1314 1178 1822 1181
rect 1826 1178 1862 1181
rect 98 1168 102 1171
rect 106 1168 286 1171
rect 426 1168 438 1171
rect 442 1168 486 1171
rect 510 1168 518 1171
rect 658 1168 686 1171
rect 690 1168 798 1171
rect 802 1168 838 1171
rect 1034 1168 1134 1171
rect 1314 1168 1502 1171
rect 1754 1168 1774 1171
rect 458 1158 502 1161
rect 510 1158 550 1161
rect 602 1158 622 1161
rect 810 1158 862 1161
rect 866 1158 1126 1161
rect 1278 1161 1281 1168
rect 1258 1158 1281 1161
rect 1362 1158 1558 1161
rect 1570 1158 1686 1161
rect 1690 1158 1726 1161
rect 1798 1158 1833 1161
rect 1842 1158 1862 1161
rect 1882 1158 1985 1161
rect 130 1148 134 1151
rect 286 1151 289 1158
rect 258 1148 289 1151
rect 354 1148 358 1151
rect 510 1151 513 1158
rect 498 1148 513 1151
rect 546 1148 582 1151
rect 602 1148 614 1151
rect 618 1148 710 1151
rect 814 1148 838 1151
rect 1074 1148 1094 1151
rect 1146 1148 1294 1151
rect 1306 1148 1310 1151
rect 1378 1148 1401 1151
rect 1426 1148 1518 1151
rect 1566 1151 1569 1158
rect 1798 1152 1801 1158
rect 1830 1152 1833 1158
rect 1982 1152 1985 1158
rect 1522 1148 1569 1151
rect 106 1138 118 1141
rect 122 1138 126 1141
rect 814 1142 817 1148
rect 1398 1142 1401 1148
rect 1650 1148 1734 1151
rect 1858 1148 1894 1151
rect 1982 1148 1986 1152
rect 146 1140 270 1141
rect 142 1138 270 1140
rect 362 1138 406 1141
rect 514 1138 630 1141
rect 866 1138 870 1141
rect 1082 1138 1206 1141
rect 1210 1138 1246 1141
rect 1298 1138 1350 1141
rect 1402 1138 1494 1141
rect 1542 1138 1742 1141
rect 1830 1141 1833 1148
rect 1830 1138 1886 1141
rect 1542 1132 1545 1138
rect 194 1128 318 1131
rect 322 1128 393 1131
rect 570 1128 606 1131
rect 778 1128 910 1131
rect 914 1128 934 1131
rect 938 1128 982 1131
rect 1106 1128 1134 1131
rect 1674 1128 1694 1131
rect 1698 1128 1766 1131
rect 1770 1128 1806 1131
rect 1858 1128 1902 1131
rect 1906 1128 1942 1131
rect 390 1122 393 1128
rect 578 1118 662 1121
rect 674 1118 854 1121
rect 1018 1118 1102 1121
rect 1234 1118 1238 1121
rect 1530 1118 1646 1121
rect 258 1108 510 1111
rect 626 1108 678 1111
rect 802 1108 894 1111
rect 898 1108 950 1111
rect 1130 1108 1230 1111
rect 1266 1108 1718 1111
rect 968 1103 970 1107
rect 974 1103 977 1107
rect 982 1103 984 1107
rect 386 1098 398 1101
rect 610 1098 766 1101
rect 874 1098 902 1101
rect 906 1098 942 1101
rect 1218 1098 1374 1101
rect 1466 1098 1470 1101
rect 1474 1098 1590 1101
rect 1594 1098 1622 1101
rect 114 1088 158 1091
rect 242 1088 270 1091
rect 370 1088 374 1091
rect 666 1088 822 1091
rect 826 1088 870 1091
rect 898 1088 918 1091
rect 954 1088 1030 1091
rect 1250 1088 1334 1091
rect 1338 1088 1358 1091
rect 1362 1088 1422 1091
rect 1426 1088 1454 1091
rect 1922 1088 1942 1091
rect 82 1078 86 1081
rect 90 1078 126 1081
rect 154 1078 166 1081
rect 298 1078 374 1081
rect 378 1078 398 1081
rect 402 1078 406 1081
rect 618 1078 638 1081
rect 650 1078 702 1081
rect 778 1078 926 1081
rect 1550 1081 1553 1088
rect 1550 1078 1606 1081
rect 1634 1078 1670 1081
rect 18 1068 78 1071
rect 82 1068 110 1071
rect 174 1071 177 1078
rect 130 1068 177 1071
rect 242 1068 305 1071
rect 370 1068 374 1071
rect 418 1068 430 1071
rect 506 1068 550 1071
rect 554 1068 654 1071
rect 658 1068 670 1071
rect 1022 1071 1025 1078
rect 1022 1068 1166 1071
rect 1382 1071 1385 1078
rect 1354 1068 1385 1071
rect 1626 1068 1646 1071
rect 1682 1068 1686 1071
rect 302 1062 305 1068
rect 590 1062 593 1068
rect 106 1058 134 1061
rect 322 1058 350 1061
rect 482 1058 486 1061
rect 650 1058 662 1061
rect 682 1058 686 1061
rect 690 1058 750 1061
rect 818 1058 838 1061
rect 898 1058 990 1061
rect 1102 1058 1134 1061
rect 1306 1058 1414 1061
rect 1526 1061 1529 1068
rect 1902 1062 1905 1068
rect 1498 1058 1529 1061
rect 1570 1058 1582 1061
rect 1610 1058 1630 1061
rect 1634 1058 1654 1061
rect 1738 1058 1822 1061
rect 1102 1052 1105 1058
rect 130 1048 142 1051
rect 202 1048 222 1051
rect 390 1048 406 1051
rect 602 1048 702 1051
rect 1226 1048 1390 1051
rect 1394 1048 1750 1051
rect 390 1042 393 1048
rect 26 1038 54 1041
rect 58 1038 190 1041
rect 426 1038 462 1041
rect 610 1038 734 1041
rect 1050 1038 1070 1041
rect 362 1028 774 1031
rect 154 1018 262 1021
rect 538 1018 558 1021
rect 562 1018 1030 1021
rect 1514 1018 1542 1021
rect 546 1008 734 1011
rect 456 1003 458 1007
rect 462 1003 465 1007
rect 470 1003 472 1007
rect 1480 1003 1482 1007
rect 1486 1003 1489 1007
rect 1494 1003 1496 1007
rect 650 998 822 1001
rect 826 998 990 1001
rect 994 998 1222 1001
rect 146 988 398 991
rect 1034 988 1118 991
rect 1186 988 1286 991
rect 1434 988 1534 991
rect 1810 988 1838 991
rect 322 978 542 981
rect 546 978 566 981
rect 570 978 606 981
rect 818 978 870 981
rect 1122 978 1126 981
rect 1162 978 1198 981
rect 362 968 422 971
rect 442 968 446 971
rect 450 968 534 971
rect 538 968 1318 971
rect 1338 968 1590 971
rect 18 958 22 961
rect 106 958 334 961
rect 350 961 353 968
rect 350 958 382 961
rect 410 958 558 961
rect 738 958 806 961
rect 810 958 1302 961
rect -26 951 -22 952
rect -26 948 6 951
rect 26 948 174 951
rect 194 948 278 951
rect 314 948 374 951
rect 394 948 398 951
rect 426 948 470 951
rect 474 948 518 951
rect 602 948 622 951
rect 682 948 742 951
rect 850 948 1214 951
rect 1258 948 1262 951
rect 1494 951 1497 958
rect 1494 948 1598 951
rect 1766 951 1769 958
rect 1746 948 1769 951
rect 1794 948 1862 951
rect 414 942 417 948
rect 582 942 585 948
rect 1662 942 1665 948
rect 1982 951 1986 952
rect 1946 948 1986 951
rect 82 938 86 941
rect 258 938 262 941
rect 338 938 358 941
rect 386 938 398 941
rect 434 938 454 941
rect 462 938 478 941
rect 874 938 934 941
rect 1082 938 1102 941
rect 1138 938 1174 941
rect 1290 938 1310 941
rect 1698 938 1726 941
rect 462 932 465 938
rect 82 928 126 931
rect 306 928 342 931
rect 394 928 430 931
rect 594 928 614 931
rect 686 931 689 938
rect 634 928 689 931
rect 810 928 878 931
rect 882 928 910 931
rect 914 928 1054 931
rect 1198 931 1201 938
rect 1198 928 1254 931
rect 1430 931 1433 938
rect 1258 928 1433 931
rect 82 918 86 921
rect 106 918 270 921
rect 346 918 422 921
rect 490 918 558 921
rect 562 918 814 921
rect 1154 918 1198 921
rect 1282 918 1310 921
rect 1322 918 1326 921
rect 1338 918 1398 921
rect 1722 918 1726 921
rect 1730 918 1910 921
rect 42 908 102 911
rect 122 908 158 911
rect 274 908 318 911
rect 458 908 582 911
rect 1306 908 1430 911
rect 1434 908 1678 911
rect 1922 908 1950 911
rect 968 903 970 907
rect 974 903 977 907
rect 982 903 984 907
rect 26 898 54 901
rect 138 898 366 901
rect 370 898 398 901
rect 410 898 510 901
rect 522 898 574 901
rect 1598 892 1601 898
rect 378 888 446 891
rect 454 888 574 891
rect 634 888 678 891
rect 1050 888 1070 891
rect 1074 888 1134 891
rect 1146 888 1238 891
rect 1842 888 1846 891
rect 454 882 457 888
rect 582 882 585 888
rect 330 878 350 881
rect 386 878 438 881
rect 538 878 582 881
rect 1066 878 1174 881
rect 1218 878 1270 881
rect 1274 878 1374 881
rect 1378 878 1422 881
rect 1426 878 1454 881
rect 1746 878 1758 881
rect 1762 878 1814 881
rect 18 868 62 871
rect 242 868 286 871
rect 290 868 358 871
rect 442 868 446 871
rect 450 868 478 871
rect 950 871 953 878
rect 950 868 1046 871
rect 1050 868 1110 871
rect 1194 868 1238 871
rect 1330 868 1374 871
rect 1378 868 1502 871
rect 1538 868 1577 871
rect 1642 868 1694 871
rect 1982 871 1986 872
rect 1954 868 1986 871
rect 78 858 86 861
rect 90 858 118 861
rect 306 858 422 861
rect 426 858 470 861
rect 602 858 606 861
rect 610 858 662 861
rect 686 861 689 868
rect 1574 862 1577 868
rect 686 858 790 861
rect 1090 858 1214 861
rect 1266 858 1382 861
rect 1386 858 1390 861
rect 1594 858 1606 861
rect 1610 858 1646 861
rect 1658 858 1665 861
rect 78 852 81 858
rect 1046 852 1049 858
rect 362 848 374 851
rect 378 848 417 851
rect 414 842 417 848
rect 466 848 478 851
rect 1406 851 1409 858
rect 1386 848 1409 851
rect 1662 852 1665 858
rect 1682 848 1750 851
rect 1754 848 1838 851
rect 1982 851 1986 852
rect 1866 848 1986 851
rect 430 841 433 848
rect 430 838 590 841
rect 1378 838 1398 841
rect 1690 838 1710 841
rect 258 828 862 831
rect 1650 828 1734 831
rect 1738 828 1782 831
rect 1786 828 1862 831
rect 154 818 166 821
rect 290 818 334 821
rect 338 818 502 821
rect 722 818 806 821
rect 810 818 1006 821
rect 1010 818 1198 821
rect 1626 818 1654 821
rect 1658 818 1710 821
rect 346 808 422 811
rect 986 808 1078 811
rect 456 803 458 807
rect 462 803 465 807
rect 470 803 472 807
rect 1480 803 1482 807
rect 1486 803 1489 807
rect 1494 803 1496 807
rect 106 798 118 801
rect 866 798 886 801
rect 890 798 990 801
rect 66 788 94 791
rect 386 788 390 791
rect 402 788 998 791
rect 1002 788 1142 791
rect 1178 788 1214 791
rect 834 778 862 781
rect 866 778 894 781
rect 898 778 1374 781
rect 322 768 454 771
rect 458 768 486 771
rect 658 768 782 771
rect 1666 768 1734 771
rect 1786 768 1806 771
rect 314 758 406 761
rect 434 758 510 761
rect 514 758 534 761
rect 558 761 561 768
rect 558 758 654 761
rect 786 758 814 761
rect 842 758 886 761
rect 922 758 1030 761
rect 1218 758 1270 761
rect 1650 758 1662 761
rect 1690 758 1702 761
rect 774 752 777 758
rect 58 748 70 751
rect 98 748 166 751
rect -26 741 -22 742
rect 6 741 9 748
rect 378 748 422 751
rect 482 748 566 751
rect 602 748 766 751
rect 802 748 814 751
rect 850 748 854 751
rect 882 748 926 751
rect 930 748 982 751
rect 1258 748 1262 751
rect 1594 748 1646 751
rect 1650 748 1662 751
rect 1798 751 1801 758
rect 1746 748 1801 751
rect -26 738 30 741
rect 74 738 142 741
rect 370 738 398 741
rect 402 738 430 741
rect 502 738 558 741
rect 562 738 574 741
rect 770 738 806 741
rect 810 738 862 741
rect 866 738 886 741
rect 1114 738 1166 741
rect 1226 738 1238 741
rect 1242 738 1286 741
rect 1346 738 1366 741
rect 1370 738 1374 741
rect 1466 738 1553 741
rect 502 732 505 738
rect 98 728 286 731
rect 290 728 398 731
rect 482 728 502 731
rect 522 728 534 731
rect 578 728 598 731
rect 630 731 633 738
rect 630 728 638 731
rect 738 728 785 731
rect 802 728 833 731
rect 1074 728 1094 731
rect 1098 728 1254 731
rect 1342 731 1345 738
rect 1550 732 1553 738
rect 1650 738 1670 741
rect 1854 741 1857 748
rect 1850 738 1857 741
rect 1282 728 1345 731
rect 1522 728 1529 731
rect 1630 731 1633 738
rect 1630 728 1694 731
rect 1714 728 1758 731
rect 782 722 785 728
rect 830 722 833 728
rect 1526 722 1529 728
rect 234 718 302 721
rect 650 718 702 721
rect 970 718 1086 721
rect 1090 718 1110 721
rect 1658 718 1678 721
rect 426 708 622 711
rect 634 708 862 711
rect 1642 708 1774 711
rect 968 703 970 707
rect 974 703 977 707
rect 982 703 984 707
rect 386 698 534 701
rect 538 698 630 701
rect 634 698 670 701
rect 778 698 958 701
rect 1402 698 1478 701
rect 1738 698 1926 701
rect 774 692 777 698
rect 626 688 630 691
rect 794 688 878 691
rect 890 688 942 691
rect 958 691 961 698
rect 958 688 974 691
rect 1170 688 1334 691
rect 1554 688 1662 691
rect 1842 688 1878 691
rect 1882 688 1934 691
rect 530 678 550 681
rect 554 678 638 681
rect 714 678 822 681
rect 826 678 878 681
rect 882 678 934 681
rect 1138 678 1238 681
rect 1242 678 1606 681
rect 1790 681 1793 688
rect 1698 678 1793 681
rect 182 668 270 671
rect 274 668 374 671
rect 698 668 734 671
rect 770 668 798 671
rect 946 668 1038 671
rect 1554 668 1590 671
rect 1634 668 1646 671
rect 1806 671 1809 678
rect 1666 668 1809 671
rect 1826 668 1870 671
rect 1982 671 1986 672
rect 1954 668 1986 671
rect 182 662 185 668
rect 418 658 430 661
rect 434 658 502 661
rect 542 661 545 668
rect 506 658 545 661
rect 570 658 598 661
rect 834 659 878 661
rect 830 658 878 659
rect 918 661 921 668
rect 882 658 921 661
rect 1070 662 1073 668
rect 1590 662 1593 668
rect 1354 658 1422 661
rect 1426 658 1470 661
rect 1534 658 1542 661
rect 1706 658 1710 661
rect 1746 658 1750 661
rect 1822 661 1825 668
rect 1786 658 1825 661
rect -26 651 -22 652
rect -26 648 6 651
rect 162 648 201 651
rect 290 648 334 651
rect 482 648 534 651
rect 538 648 590 651
rect 1650 648 1734 651
rect 1982 651 1986 652
rect 1914 648 1986 651
rect 198 642 201 648
rect 282 638 846 641
rect 850 638 1222 641
rect 1226 638 1246 641
rect 1602 638 1630 641
rect 1634 638 1694 641
rect 34 628 1238 631
rect 1242 628 1406 631
rect 1610 628 1622 631
rect 1626 628 1718 631
rect 186 618 222 621
rect 226 618 294 621
rect 298 618 366 621
rect 456 603 458 607
rect 462 603 465 607
rect 470 603 472 607
rect 1480 603 1482 607
rect 1486 603 1489 607
rect 1494 603 1496 607
rect 354 598 382 601
rect 1934 592 1937 598
rect 698 588 734 591
rect 514 578 806 581
rect 1402 578 1406 581
rect 1410 578 1494 581
rect 1498 578 1638 581
rect 1674 578 1694 581
rect 1698 578 1702 581
rect 98 568 129 571
rect 202 568 254 571
rect 482 568 726 571
rect 730 568 758 571
rect 1058 568 1102 571
rect 1482 568 1697 571
rect 1786 568 1854 571
rect 1858 568 1862 571
rect 126 562 129 568
rect 806 562 809 568
rect 90 558 102 561
rect 322 558 358 561
rect 378 558 398 561
rect 402 558 446 561
rect 458 558 494 561
rect 498 558 518 561
rect 522 558 614 561
rect 618 558 766 561
rect 830 558 838 561
rect 842 558 862 561
rect 874 558 1038 561
rect 1058 558 1118 561
rect 1158 561 1161 568
rect 1694 562 1697 568
rect 1122 558 1161 561
rect 1606 558 1630 561
rect 1698 558 1710 561
rect 1722 558 1798 561
rect 102 551 105 558
rect 230 551 233 558
rect 1606 552 1609 558
rect 102 548 478 551
rect 490 548 510 551
rect 578 548 670 551
rect 674 548 710 551
rect 762 548 878 551
rect 1090 548 1126 551
rect 1134 548 1142 551
rect 1178 548 1214 551
rect 1458 548 1470 551
rect 1530 548 1593 551
rect 1674 548 1758 551
rect 1778 548 1798 551
rect 1590 542 1593 548
rect 18 538 30 541
rect 114 538 142 541
rect 226 538 246 541
rect 586 538 646 541
rect 730 538 774 541
rect 842 538 846 541
rect 882 538 1086 541
rect 1090 538 1094 541
rect 1098 538 1182 541
rect 1194 538 1198 541
rect 1210 538 1302 541
rect 1682 538 1710 541
rect 1730 538 1766 541
rect 1770 538 1782 541
rect 1794 538 1822 541
rect 242 528 278 531
rect 282 528 302 531
rect 426 528 478 531
rect 578 528 726 531
rect 730 528 838 531
rect 866 528 870 531
rect 906 528 934 531
rect 1034 528 1134 531
rect 1154 528 1366 531
rect 1522 528 1558 531
rect 1618 528 1726 531
rect 1938 528 1942 531
rect 710 522 713 528
rect 842 518 982 521
rect 1146 518 1238 521
rect 1570 518 1654 521
rect 1122 508 1390 511
rect 1394 508 1598 511
rect 968 503 970 507
rect 974 503 977 507
rect 982 503 984 507
rect 186 498 214 501
rect 218 498 278 501
rect 410 498 430 501
rect 1626 498 1686 501
rect 1722 498 1806 501
rect 42 488 110 491
rect 114 488 286 491
rect 334 491 337 498
rect 306 488 337 491
rect 382 492 385 498
rect 790 492 793 498
rect 886 492 889 498
rect 394 488 430 491
rect 490 488 686 491
rect 998 488 1006 491
rect 1010 488 1190 491
rect 1194 488 1374 491
rect 1402 488 1526 491
rect 1594 488 1646 491
rect 1650 488 1806 491
rect 1810 488 1838 491
rect 90 478 134 481
rect 138 478 158 481
rect 306 478 558 481
rect 682 478 686 481
rect 810 478 830 481
rect 834 478 902 481
rect 906 478 1062 481
rect 1442 478 1513 481
rect 1538 478 1694 481
rect 330 468 374 471
rect 558 471 561 478
rect 558 468 582 471
rect 638 471 641 478
rect 1510 472 1513 478
rect 638 468 646 471
rect 826 468 918 471
rect 922 468 1046 471
rect 1050 468 1070 471
rect 1074 468 1198 471
rect 1202 468 1246 471
rect 1266 468 1302 471
rect 1306 468 1350 471
rect 1690 468 1694 471
rect 538 459 742 461
rect 534 458 742 459
rect 906 458 926 461
rect 930 458 950 461
rect 1018 458 1150 461
rect 1454 461 1457 468
rect 1338 458 1526 461
rect 1554 458 1558 461
rect 1578 458 1582 461
rect 1642 459 1710 461
rect 1638 458 1710 459
rect 1750 461 1753 468
rect 1854 462 1857 468
rect 1714 458 1753 461
rect 1802 458 1846 461
rect -26 451 -22 452
rect -26 448 6 451
rect 914 448 990 451
rect 1162 448 1686 451
rect 850 438 1102 441
rect 1570 438 1614 441
rect 1618 438 1662 441
rect 362 428 374 431
rect 1554 428 1574 431
rect 1578 428 1710 431
rect 1714 428 1782 431
rect 456 403 458 407
rect 462 403 465 407
rect 470 403 472 407
rect 1480 403 1482 407
rect 1486 403 1489 407
rect 1494 403 1496 407
rect 98 398 222 401
rect 18 388 78 391
rect 82 388 94 391
rect 410 388 526 391
rect 890 388 958 391
rect 962 388 974 391
rect 978 388 1062 391
rect 1122 368 1182 371
rect 1186 368 1214 371
rect 290 358 390 361
rect 482 358 502 361
rect 70 351 73 358
rect 70 348 142 351
rect 402 348 406 351
rect 458 348 518 351
rect 694 351 697 358
rect 682 348 697 351
rect 918 351 921 358
rect 858 348 921 351
rect 1190 351 1193 358
rect 1238 352 1241 358
rect 1190 348 1206 351
rect 1522 348 1622 351
rect 1678 348 1686 351
rect 1690 348 1742 351
rect 1746 348 1750 351
rect 250 338 326 341
rect 362 338 422 341
rect 498 338 510 341
rect 730 338 750 341
rect 754 338 990 341
rect 994 340 1014 341
rect 1390 342 1393 348
rect 994 338 1017 340
rect 1042 338 1054 341
rect 1058 338 1134 341
rect 1450 338 1734 341
rect 1582 332 1585 338
rect 506 328 534 331
rect 654 328 678 331
rect 794 328 838 331
rect 954 328 1038 331
rect 1042 328 1126 331
rect 654 322 657 328
rect 306 318 398 321
rect 386 308 430 311
rect 1090 308 1206 311
rect 1210 308 1238 311
rect 1242 308 1294 311
rect 1298 308 1350 311
rect 968 303 970 307
rect 974 303 977 307
rect 982 303 984 307
rect 66 298 110 301
rect 1682 298 1702 301
rect 354 288 369 291
rect 402 288 478 291
rect 1554 288 1622 291
rect 1658 288 1670 291
rect 1794 288 1822 291
rect 366 282 369 288
rect 686 281 689 288
rect 686 278 766 281
rect 1674 278 1686 281
rect 1774 281 1777 288
rect 1690 278 1777 281
rect 286 271 289 278
rect 406 271 409 278
rect 146 268 409 271
rect 958 271 961 278
rect 922 268 1054 271
rect 1290 268 1390 271
rect 130 258 209 261
rect 386 258 398 261
rect 754 258 774 261
rect 1242 258 1337 261
rect 1498 258 1577 261
rect 1602 258 1718 261
rect 1722 258 1806 261
rect 126 252 129 258
rect 206 252 209 258
rect -26 251 -22 252
rect -26 248 6 251
rect 10 248 38 251
rect 42 248 70 251
rect 682 248 694 251
rect 1238 251 1241 258
rect 698 248 1241 251
rect 1334 252 1337 258
rect 1574 252 1577 258
rect 82 238 510 241
rect 514 238 734 241
rect 762 238 782 241
rect 818 238 1374 241
rect 1378 238 1454 241
rect 258 228 302 231
rect 306 228 406 231
rect 722 228 742 231
rect 186 218 262 221
rect 794 218 806 221
rect 810 218 870 221
rect 922 218 1486 221
rect 1026 208 1118 211
rect 456 203 458 207
rect 462 203 465 207
rect 470 203 472 207
rect 1480 203 1482 207
rect 1486 203 1489 207
rect 1494 203 1496 207
rect 1090 198 1110 201
rect 1114 198 1174 201
rect 850 188 934 191
rect 1434 188 1518 191
rect 1738 188 1774 191
rect 878 182 881 188
rect 210 168 238 171
rect 474 168 486 171
rect 758 171 761 178
rect 698 168 761 171
rect 114 158 414 161
rect 602 158 670 161
rect 754 158 774 161
rect 794 158 814 161
rect 1346 158 1398 161
rect 1402 158 1542 161
rect 1770 158 1798 161
rect 1802 158 1886 161
rect -26 151 -22 152
rect -26 148 6 151
rect 90 148 177 151
rect 194 148 238 151
rect 298 148 318 151
rect 322 148 350 151
rect 562 148 886 151
rect 890 148 1094 151
rect 1098 148 1102 151
rect 1106 148 1254 151
rect 1278 151 1281 158
rect 1278 148 1318 151
rect 1418 148 1438 151
rect 1554 148 1558 151
rect 1690 148 1726 151
rect 1842 148 1878 151
rect 174 142 177 148
rect 574 138 598 141
rect 650 138 654 141
rect 818 138 838 141
rect 874 138 918 141
rect 1010 138 1078 141
rect 1082 138 1142 141
rect 1194 138 1310 141
rect 1366 141 1369 148
rect 1314 138 1369 141
rect 1394 138 1422 141
rect 1554 138 1646 141
rect 1650 138 1694 141
rect 1698 138 1782 141
rect 1834 138 1838 141
rect 262 131 265 138
rect 286 131 289 138
rect 574 132 577 138
rect 262 128 289 131
rect 434 128 574 131
rect 618 128 782 131
rect 786 128 822 131
rect 826 128 926 131
rect 930 128 1542 131
rect 1546 128 1814 131
rect 1830 128 1942 131
rect 1830 122 1833 128
rect 10 118 38 121
rect 42 118 142 121
rect 146 118 230 121
rect 234 118 270 121
rect 274 118 302 121
rect 418 118 502 121
rect 506 118 550 121
rect 794 118 814 121
rect 826 118 902 121
rect 906 118 990 121
rect 1010 118 1046 121
rect 1050 118 1057 121
rect 1210 118 1358 121
rect 1362 118 1406 121
rect 1586 118 1622 121
rect 1674 118 1702 121
rect 1706 118 1726 121
rect 1778 118 1806 121
rect 1810 118 1830 121
rect 74 108 134 111
rect 306 108 454 111
rect 458 108 462 111
rect 642 108 790 111
rect 802 108 822 111
rect 1042 108 1054 111
rect 1066 108 1150 111
rect 1154 108 1398 111
rect 968 103 970 107
rect 974 103 977 107
rect 982 103 984 107
rect 122 98 126 101
rect 130 98 270 101
rect 418 98 622 101
rect 626 98 670 101
rect 818 98 862 101
rect 1162 98 1206 101
rect 1354 98 1369 101
rect 1378 98 1390 101
rect 1394 98 1502 101
rect 1366 92 1369 98
rect 118 88 126 91
rect 218 88 310 91
rect 362 88 470 91
rect 794 88 862 91
rect 1010 88 1038 91
rect 1234 88 1262 91
rect 1266 88 1366 91
rect 1418 88 1446 91
rect 1450 88 1582 91
rect 1626 88 1670 91
rect 1674 88 1758 91
rect 130 78 134 81
rect 170 78 206 81
rect 242 78 294 81
rect 298 78 326 81
rect 338 78 486 81
rect 606 81 609 88
rect 490 78 609 81
rect 750 81 753 88
rect 918 82 921 88
rect 750 78 798 81
rect 930 78 1150 81
rect 1214 81 1217 88
rect 1154 78 1217 81
rect 1234 78 1246 81
rect 1298 78 1454 81
rect 1634 78 1718 81
rect 1722 78 1782 81
rect 114 68 118 71
rect 162 68 174 71
rect 178 68 230 71
rect 346 68 518 71
rect 522 68 590 71
rect 594 68 614 71
rect 778 68 790 71
rect 858 68 878 71
rect 886 71 889 78
rect 882 68 889 71
rect 894 68 998 71
rect 1010 68 1014 71
rect 1026 68 1030 71
rect 1074 68 1118 71
rect 1294 71 1297 78
rect 1138 68 1297 71
rect 1594 68 1758 71
rect 1854 71 1857 78
rect 1762 68 1857 71
rect 42 58 150 61
rect 154 58 161 61
rect 170 58 598 61
rect 602 58 638 61
rect 894 61 897 68
rect 642 58 897 61
rect 986 58 1046 61
rect 1050 58 1086 61
rect 1090 58 1198 61
rect 1202 58 1233 61
rect 1242 58 1270 61
rect 1282 58 1390 61
rect 1578 58 1630 61
rect 1634 58 1678 61
rect 1786 58 1825 61
rect 1230 52 1233 58
rect 1822 52 1825 58
rect 50 48 54 51
rect 146 48 158 51
rect 178 48 198 51
rect 202 48 334 51
rect 418 48 422 51
rect 498 48 510 51
rect 522 48 550 51
rect 858 48 878 51
rect 882 48 1182 51
rect 1186 48 1222 51
rect 1266 48 1334 51
rect 258 38 294 41
rect 298 38 534 41
rect 538 38 846 41
rect 1034 38 1070 41
rect 1222 41 1225 48
rect 1222 38 1630 41
rect 766 22 769 28
rect 456 3 458 7
rect 462 3 465 7
rect 470 3 472 7
rect 1480 3 1482 7
rect 1486 3 1489 7
rect 1494 3 1496 7
<< m4contact >>
rect 970 1703 974 1707
rect 978 1703 981 1707
rect 981 1703 982 1707
rect 1070 1698 1074 1702
rect 1150 1698 1154 1702
rect 1318 1698 1322 1702
rect 1158 1658 1162 1662
rect 1022 1638 1026 1642
rect 1326 1628 1330 1632
rect 862 1618 866 1622
rect 1246 1618 1250 1622
rect 1654 1618 1658 1622
rect 1062 1608 1066 1612
rect 458 1603 462 1607
rect 466 1603 469 1607
rect 469 1603 470 1607
rect 1482 1603 1486 1607
rect 1490 1603 1493 1607
rect 1493 1603 1494 1607
rect 438 1578 442 1582
rect 1742 1548 1746 1552
rect 606 1538 610 1542
rect 958 1528 962 1532
rect 1654 1528 1658 1532
rect 814 1508 818 1512
rect 970 1503 974 1507
rect 978 1503 981 1507
rect 981 1503 982 1507
rect 1022 1478 1026 1482
rect 1230 1478 1234 1482
rect 1622 1478 1626 1482
rect 406 1468 410 1472
rect 1230 1458 1234 1462
rect 958 1448 962 1452
rect 1246 1448 1250 1452
rect 1622 1448 1626 1452
rect 126 1438 130 1442
rect 1222 1438 1226 1442
rect 1382 1428 1386 1432
rect 1902 1428 1906 1432
rect 458 1403 462 1407
rect 466 1403 469 1407
rect 469 1403 470 1407
rect 1482 1403 1486 1407
rect 1490 1403 1493 1407
rect 1493 1403 1494 1407
rect 446 1388 450 1392
rect 1590 1388 1594 1392
rect 790 1378 794 1382
rect 1118 1378 1122 1382
rect 1734 1378 1738 1382
rect 734 1368 738 1372
rect 278 1358 282 1362
rect 374 1358 378 1362
rect 118 1348 122 1352
rect 758 1348 762 1352
rect 926 1348 930 1352
rect 1230 1348 1234 1352
rect 1302 1348 1306 1352
rect 1654 1348 1658 1352
rect 566 1338 570 1342
rect 1414 1338 1418 1342
rect 1582 1338 1586 1342
rect 758 1328 762 1332
rect 894 1308 898 1312
rect 970 1303 974 1307
rect 978 1303 981 1307
rect 981 1303 982 1307
rect 846 1298 850 1302
rect 806 1278 810 1282
rect 270 1268 274 1272
rect 1222 1268 1226 1272
rect 1598 1268 1602 1272
rect 1934 1268 1938 1272
rect 150 1258 154 1262
rect 598 1258 602 1262
rect 382 1248 386 1252
rect 406 1248 410 1252
rect 734 1248 738 1252
rect 1398 1248 1402 1252
rect 598 1238 602 1242
rect 1382 1238 1386 1242
rect 1654 1238 1658 1242
rect 574 1228 578 1232
rect 1286 1228 1290 1232
rect 1742 1218 1746 1222
rect 478 1208 482 1212
rect 458 1203 462 1207
rect 466 1203 469 1207
rect 469 1203 470 1207
rect 1482 1203 1486 1207
rect 1490 1203 1493 1207
rect 1493 1203 1494 1207
rect 822 1198 826 1202
rect 1398 1188 1402 1192
rect 94 1168 98 1172
rect 358 1148 362 1152
rect 598 1148 602 1152
rect 1302 1148 1306 1152
rect 126 1138 130 1142
rect 270 1138 274 1142
rect 870 1138 874 1142
rect 1942 1128 1946 1132
rect 1230 1118 1234 1122
rect 798 1108 802 1112
rect 970 1103 974 1107
rect 978 1103 981 1107
rect 981 1103 982 1107
rect 606 1098 610 1102
rect 270 1088 274 1092
rect 374 1088 378 1092
rect 398 1078 402 1082
rect 926 1078 930 1082
rect 126 1068 130 1072
rect 374 1068 378 1072
rect 502 1068 506 1072
rect 486 1058 490 1062
rect 814 1058 818 1062
rect 1734 1058 1738 1062
rect 1902 1058 1906 1062
rect 1390 1048 1394 1052
rect 358 1028 362 1032
rect 558 1018 562 1022
rect 458 1003 462 1007
rect 466 1003 469 1007
rect 469 1003 470 1007
rect 1482 1003 1486 1007
rect 1490 1003 1493 1007
rect 1493 1003 1494 1007
rect 646 998 650 1002
rect 1286 988 1290 992
rect 1126 978 1130 982
rect 422 968 426 972
rect 438 968 442 972
rect 102 958 106 962
rect 406 958 410 962
rect 1302 958 1306 962
rect 174 948 178 952
rect 398 948 402 952
rect 414 948 418 952
rect 422 948 426 952
rect 1262 948 1266 952
rect 1662 948 1666 952
rect 86 938 90 942
rect 254 938 258 942
rect 454 938 458 942
rect 582 938 586 942
rect 1286 938 1290 942
rect 78 918 82 922
rect 1326 918 1330 922
rect 102 908 106 912
rect 158 908 162 912
rect 454 908 458 912
rect 1302 908 1306 912
rect 970 903 974 907
rect 978 903 981 907
rect 981 903 982 907
rect 398 898 402 902
rect 510 898 514 902
rect 374 888 378 892
rect 574 888 578 892
rect 1046 888 1050 892
rect 1598 888 1602 892
rect 1846 888 1850 892
rect 582 878 586 882
rect 438 868 442 872
rect 86 858 90 862
rect 118 858 122 862
rect 598 858 602 862
rect 1046 858 1050 862
rect 1382 858 1386 862
rect 1646 858 1650 862
rect 478 848 482 852
rect 1862 848 1866 852
rect 1398 838 1402 842
rect 502 818 506 822
rect 806 818 810 822
rect 1710 818 1714 822
rect 458 803 462 807
rect 466 803 469 807
rect 469 803 470 807
rect 1482 803 1486 807
rect 1490 803 1493 807
rect 1493 803 1494 807
rect 886 798 890 802
rect 382 788 386 792
rect 398 788 402 792
rect 894 778 898 782
rect 406 758 410 762
rect 782 758 786 762
rect 774 748 778 752
rect 798 748 802 752
rect 846 748 850 752
rect 1254 748 1258 752
rect 1662 748 1666 752
rect 398 738 402 742
rect 1222 738 1226 742
rect 638 728 642 732
rect 1070 728 1074 732
rect 1846 738 1850 742
rect 1518 728 1522 732
rect 1710 728 1714 732
rect 630 708 634 712
rect 970 703 974 707
rect 978 703 981 707
rect 981 703 982 707
rect 630 688 634 692
rect 774 688 778 692
rect 1238 678 1242 682
rect 798 668 802 672
rect 1070 658 1074 662
rect 1590 658 1594 662
rect 1710 658 1714 662
rect 478 648 482 652
rect 846 638 850 642
rect 458 603 462 607
rect 466 603 469 607
rect 469 603 470 607
rect 1482 603 1486 607
rect 1490 603 1493 607
rect 1493 603 1494 607
rect 1934 588 1938 592
rect 806 578 810 582
rect 1694 578 1698 582
rect 478 568 482 572
rect 806 568 810 572
rect 1854 568 1858 572
rect 86 558 90 562
rect 478 548 482 552
rect 1142 548 1146 552
rect 846 538 850 542
rect 1190 538 1194 542
rect 1782 538 1786 542
rect 1942 528 1946 532
rect 838 518 842 522
rect 970 503 974 507
rect 978 503 981 507
rect 981 503 982 507
rect 790 498 794 502
rect 382 488 386 492
rect 886 488 890 492
rect 1838 488 1842 492
rect 678 478 682 482
rect 646 468 650 472
rect 1694 468 1698 472
rect 1854 458 1858 462
rect 374 428 378 432
rect 1710 428 1714 432
rect 458 403 462 407
rect 466 403 469 407
rect 469 403 470 407
rect 1482 403 1486 407
rect 1490 403 1493 407
rect 1493 403 1494 407
rect 78 388 82 392
rect 398 348 402 352
rect 1238 348 1242 352
rect 1390 338 1394 342
rect 838 328 842 332
rect 398 318 402 322
rect 970 303 974 307
rect 978 303 981 307
rect 981 303 982 307
rect 398 288 402 292
rect 766 278 770 282
rect 918 268 922 272
rect 398 258 402 262
rect 1238 258 1242 262
rect 126 248 130 252
rect 678 248 682 252
rect 458 203 462 207
rect 466 203 469 207
rect 469 203 470 207
rect 1482 203 1486 207
rect 1490 203 1493 207
rect 1493 203 1494 207
rect 1518 188 1522 192
rect 790 158 794 162
rect 1558 148 1562 152
rect 654 138 658 142
rect 1142 138 1146 142
rect 1830 138 1834 142
rect 414 118 418 122
rect 790 108 794 112
rect 970 103 974 107
rect 978 103 981 107
rect 981 103 982 107
rect 118 98 122 102
rect 126 88 130 92
rect 126 78 130 82
rect 334 78 338 82
rect 886 78 890 82
rect 918 78 922 82
rect 118 68 122 72
rect 1014 68 1018 72
rect 1030 68 1034 72
rect 1238 58 1242 62
rect 1782 58 1786 62
rect 46 48 50 52
rect 174 48 178 52
rect 334 48 338 52
rect 422 48 426 52
rect 518 48 522 52
rect 766 28 770 32
rect 458 3 462 7
rect 466 3 469 7
rect 469 3 470 7
rect 1482 3 1486 7
rect 1490 3 1493 7
rect 1493 3 1494 7
<< metal4 >>
rect 968 1703 970 1707
rect 974 1703 977 1707
rect 982 1703 984 1707
rect 1062 1698 1070 1701
rect 1154 1698 1161 1701
rect 1322 1698 1329 1701
rect 456 1603 458 1607
rect 462 1603 465 1607
rect 470 1603 472 1607
rect 442 1578 449 1581
rect 98 1168 105 1171
rect 102 962 105 1168
rect 78 938 86 941
rect 78 922 81 938
rect 78 392 81 918
rect 102 912 105 958
rect 118 862 121 1348
rect 126 1142 129 1438
rect 270 1358 278 1361
rect 270 1272 273 1358
rect 154 1258 161 1261
rect 126 1072 129 1138
rect 158 912 161 1258
rect 270 1142 273 1268
rect 374 1251 377 1358
rect 406 1252 409 1468
rect 446 1392 449 1578
rect 456 1403 458 1407
rect 462 1403 465 1407
rect 470 1403 472 1407
rect 558 1338 566 1341
rect 374 1248 382 1251
rect 270 1092 273 1138
rect 358 1032 361 1148
rect 374 1072 377 1088
rect 406 1081 409 1248
rect 456 1203 458 1207
rect 462 1203 465 1207
rect 470 1203 472 1207
rect 402 1078 409 1081
rect 478 1061 481 1208
rect 478 1058 486 1061
rect 456 1003 458 1007
rect 462 1003 465 1007
rect 470 1003 472 1007
rect 178 948 182 951
rect 394 948 398 951
rect 258 938 262 941
rect 86 562 89 858
rect 374 432 377 888
rect 398 792 401 898
rect 382 492 385 788
rect 406 762 409 958
rect 422 952 425 968
rect 414 942 417 948
rect 438 872 441 968
rect 454 912 457 938
rect 456 803 458 807
rect 462 803 465 807
rect 470 803 472 807
rect 398 352 401 738
rect 478 652 481 848
rect 502 822 505 1068
rect 558 1022 561 1338
rect 598 1242 601 1258
rect 510 902 513 918
rect 574 892 577 1228
rect 582 882 585 938
rect 598 862 601 1148
rect 606 1102 609 1538
rect 806 1508 814 1511
rect 734 1252 737 1368
rect 758 1332 761 1348
rect 638 732 641 738
rect 630 692 633 708
rect 456 603 458 607
rect 462 603 465 607
rect 470 603 472 607
rect 478 552 481 568
rect 646 472 649 998
rect 774 692 777 748
rect 782 732 785 758
rect 790 502 793 1378
rect 806 1282 809 1508
rect 814 1198 822 1201
rect 798 752 801 1108
rect 814 1062 817 1198
rect 798 672 801 748
rect 806 582 809 818
rect 846 752 849 1298
rect 862 1141 865 1618
rect 958 1452 961 1528
rect 968 1503 970 1507
rect 974 1503 977 1507
rect 982 1503 984 1507
rect 1022 1482 1025 1638
rect 1062 1612 1065 1698
rect 1158 1662 1161 1698
rect 1326 1632 1329 1698
rect 1230 1462 1233 1478
rect 1246 1452 1249 1618
rect 1480 1603 1482 1607
rect 1486 1603 1489 1607
rect 1494 1603 1496 1607
rect 1654 1532 1657 1618
rect 1622 1452 1625 1478
rect 862 1138 870 1141
rect 846 642 849 748
rect 806 572 809 578
rect 838 538 846 541
rect 838 522 841 538
rect 456 403 458 407
rect 462 403 465 407
rect 470 403 472 407
rect 398 322 401 348
rect 398 292 401 318
rect 398 262 401 288
rect 118 72 121 98
rect 126 92 129 248
rect 456 203 458 207
rect 462 203 465 207
rect 470 203 472 207
rect 646 141 649 468
rect 678 252 681 478
rect 838 332 841 518
rect 886 492 889 798
rect 894 782 897 1308
rect 926 1082 929 1348
rect 968 1303 970 1307
rect 974 1303 977 1307
rect 982 1303 984 1307
rect 968 1103 970 1107
rect 974 1103 977 1107
rect 982 1103 984 1107
rect 1118 981 1121 1378
rect 1222 1272 1225 1438
rect 1118 978 1126 981
rect 968 903 970 907
rect 974 903 977 907
rect 982 903 984 907
rect 1046 862 1049 888
rect 1222 742 1225 1268
rect 1230 1122 1233 1348
rect 1286 992 1289 1228
rect 1302 1152 1305 1348
rect 1382 1242 1385 1428
rect 1480 1403 1482 1407
rect 1486 1403 1489 1407
rect 1494 1403 1496 1407
rect 1418 1338 1422 1341
rect 1578 1338 1582 1341
rect 1254 948 1262 951
rect 1254 752 1257 948
rect 1286 942 1289 988
rect 1302 962 1305 1148
rect 1302 912 1305 958
rect 1322 918 1326 921
rect 1382 862 1385 1238
rect 1398 1192 1401 1248
rect 1480 1203 1482 1207
rect 1486 1203 1489 1207
rect 1494 1203 1496 1207
rect 968 703 970 707
rect 974 703 977 707
rect 982 703 984 707
rect 1070 662 1073 728
rect 1142 542 1145 548
rect 1194 538 1198 541
rect 968 503 970 507
rect 974 503 977 507
rect 982 503 984 507
rect 1238 352 1241 678
rect 968 303 970 307
rect 974 303 977 307
rect 982 303 984 307
rect 646 138 654 141
rect 130 78 134 81
rect 334 52 337 78
rect 50 48 54 51
rect 170 48 174 51
rect 414 51 417 118
rect 518 52 521 78
rect 414 48 422 51
rect 766 32 769 278
rect 790 112 793 158
rect 918 82 921 268
rect 1238 262 1241 348
rect 1390 342 1393 1048
rect 1398 842 1401 1188
rect 1480 1003 1482 1007
rect 1486 1003 1489 1007
rect 1494 1003 1496 1007
rect 1480 803 1482 807
rect 1486 803 1489 807
rect 1494 803 1496 807
rect 1480 603 1482 607
rect 1486 603 1489 607
rect 1494 603 1496 607
rect 1480 403 1482 407
rect 1486 403 1489 407
rect 1494 403 1496 407
rect 1480 203 1482 207
rect 1486 203 1489 207
rect 1494 203 1496 207
rect 1518 192 1521 728
rect 1590 662 1593 1388
rect 1654 1352 1657 1528
rect 1598 892 1601 1268
rect 1654 1242 1657 1348
rect 1734 1062 1737 1378
rect 1742 1222 1745 1548
rect 1902 1062 1905 1428
rect 1646 852 1649 858
rect 1662 752 1665 948
rect 1710 732 1713 818
rect 1846 742 1849 888
rect 1858 848 1862 851
rect 1710 662 1713 728
rect 1694 472 1697 578
rect 1710 432 1713 658
rect 1934 592 1937 1268
rect 1554 148 1558 151
rect 1142 142 1145 148
rect 968 103 970 107
rect 974 103 977 107
rect 982 103 984 107
rect 886 72 889 78
rect 1010 68 1014 71
rect 1026 68 1030 71
rect 1238 62 1241 68
rect 1782 62 1785 538
rect 1838 141 1841 488
rect 1854 462 1857 568
rect 1942 532 1945 1128
rect 1834 138 1841 141
rect 456 3 458 7
rect 462 3 465 7
rect 470 3 472 7
rect 1480 3 1482 7
rect 1486 3 1489 7
rect 1494 3 1496 7
<< m5contact >>
rect 970 1703 974 1707
rect 977 1703 978 1707
rect 978 1703 981 1707
rect 458 1603 462 1607
rect 465 1603 466 1607
rect 466 1603 469 1607
rect 458 1403 462 1407
rect 465 1403 466 1407
rect 466 1403 469 1407
rect 458 1203 462 1207
rect 465 1203 466 1207
rect 466 1203 469 1207
rect 458 1003 462 1007
rect 465 1003 466 1007
rect 466 1003 469 1007
rect 182 948 186 952
rect 390 948 394 952
rect 262 938 266 942
rect 414 938 418 942
rect 458 803 462 807
rect 465 803 466 807
rect 466 803 469 807
rect 510 918 514 922
rect 638 738 642 742
rect 458 603 462 607
rect 465 603 466 607
rect 466 603 469 607
rect 782 728 786 732
rect 970 1503 974 1507
rect 977 1503 978 1507
rect 978 1503 981 1507
rect 1482 1603 1486 1607
rect 1489 1603 1490 1607
rect 1490 1603 1493 1607
rect 458 403 462 407
rect 465 403 466 407
rect 466 403 469 407
rect 458 203 462 207
rect 465 203 466 207
rect 466 203 469 207
rect 970 1303 974 1307
rect 977 1303 978 1307
rect 978 1303 981 1307
rect 970 1103 974 1107
rect 977 1103 978 1107
rect 978 1103 981 1107
rect 970 903 974 907
rect 977 903 978 907
rect 978 903 981 907
rect 1482 1403 1486 1407
rect 1489 1403 1490 1407
rect 1490 1403 1493 1407
rect 1422 1338 1426 1342
rect 1574 1338 1578 1342
rect 1318 918 1322 922
rect 1482 1203 1486 1207
rect 1489 1203 1490 1207
rect 1490 1203 1493 1207
rect 970 703 974 707
rect 977 703 978 707
rect 978 703 981 707
rect 1142 538 1146 542
rect 1198 538 1202 542
rect 970 503 974 507
rect 977 503 978 507
rect 978 503 981 507
rect 970 303 974 307
rect 977 303 978 307
rect 978 303 981 307
rect 134 78 138 82
rect 54 48 58 52
rect 166 48 170 52
rect 518 78 522 82
rect 1482 1003 1486 1007
rect 1489 1003 1490 1007
rect 1490 1003 1493 1007
rect 1482 803 1486 807
rect 1489 803 1490 807
rect 1490 803 1493 807
rect 1482 603 1486 607
rect 1489 603 1490 607
rect 1490 603 1493 607
rect 1482 403 1486 407
rect 1489 403 1490 407
rect 1490 403 1493 407
rect 1482 203 1486 207
rect 1489 203 1490 207
rect 1490 203 1493 207
rect 1646 848 1650 852
rect 1854 848 1858 852
rect 1142 148 1146 152
rect 1550 148 1554 152
rect 970 103 974 107
rect 977 103 978 107
rect 978 103 981 107
rect 886 68 890 72
rect 1006 68 1010 72
rect 1022 68 1026 72
rect 1238 68 1242 72
rect 458 3 462 7
rect 465 3 466 7
rect 466 3 469 7
rect 1482 3 1486 7
rect 1489 3 1490 7
rect 1490 3 1493 7
<< metal5 >>
rect 974 1703 977 1707
rect 973 1702 978 1703
rect 983 1702 984 1707
rect 462 1603 465 1607
rect 461 1602 466 1603
rect 471 1602 472 1607
rect 1486 1603 1489 1607
rect 1485 1602 1490 1603
rect 1495 1602 1496 1607
rect 974 1503 977 1507
rect 973 1502 978 1503
rect 983 1502 984 1507
rect 462 1403 465 1407
rect 461 1402 466 1403
rect 471 1402 472 1407
rect 1486 1403 1489 1407
rect 1485 1402 1490 1403
rect 1495 1402 1496 1407
rect 1426 1338 1574 1341
rect 974 1303 977 1307
rect 973 1302 978 1303
rect 983 1302 984 1307
rect 462 1203 465 1207
rect 461 1202 466 1203
rect 471 1202 472 1207
rect 1486 1203 1489 1207
rect 1485 1202 1490 1203
rect 1495 1202 1496 1207
rect 974 1103 977 1107
rect 973 1102 978 1103
rect 983 1102 984 1107
rect 462 1003 465 1007
rect 461 1002 466 1003
rect 471 1002 472 1007
rect 1486 1003 1489 1007
rect 1485 1002 1490 1003
rect 1495 1002 1496 1007
rect 186 948 390 951
rect 266 938 414 941
rect 514 918 1318 921
rect 974 903 977 907
rect 973 902 978 903
rect 983 902 984 907
rect 1650 848 1854 851
rect 462 803 465 807
rect 461 802 466 803
rect 471 802 472 807
rect 1486 803 1489 807
rect 1485 802 1490 803
rect 1495 802 1496 807
rect 638 731 641 738
rect 638 728 782 731
rect 974 703 977 707
rect 973 702 978 703
rect 983 702 984 707
rect 462 603 465 607
rect 461 602 466 603
rect 471 602 472 607
rect 1486 603 1489 607
rect 1485 602 1490 603
rect 1495 602 1496 607
rect 1146 538 1198 541
rect 974 503 977 507
rect 973 502 978 503
rect 983 502 984 507
rect 462 403 465 407
rect 461 402 466 403
rect 471 402 472 407
rect 1486 403 1489 407
rect 1485 402 1490 403
rect 1495 402 1496 407
rect 974 303 977 307
rect 973 302 978 303
rect 983 302 984 307
rect 462 203 465 207
rect 461 202 466 203
rect 471 202 472 207
rect 1486 203 1489 207
rect 1485 202 1490 203
rect 1495 202 1496 207
rect 1146 148 1550 151
rect 974 103 977 107
rect 973 102 978 103
rect 983 102 984 107
rect 138 78 518 81
rect 890 68 1006 71
rect 1026 68 1238 71
rect 58 48 166 51
rect 462 3 465 7
rect 461 2 466 3
rect 471 2 472 7
rect 1486 3 1489 7
rect 1485 2 1490 3
rect 1495 2 1496 7
<< m6contact >>
rect 968 1703 970 1707
rect 970 1703 973 1707
rect 978 1703 981 1707
rect 981 1703 983 1707
rect 968 1702 973 1703
rect 978 1702 983 1703
rect 456 1603 458 1607
rect 458 1603 461 1607
rect 466 1603 469 1607
rect 469 1603 471 1607
rect 456 1602 461 1603
rect 466 1602 471 1603
rect 1480 1603 1482 1607
rect 1482 1603 1485 1607
rect 1490 1603 1493 1607
rect 1493 1603 1495 1607
rect 1480 1602 1485 1603
rect 1490 1602 1495 1603
rect 968 1503 970 1507
rect 970 1503 973 1507
rect 978 1503 981 1507
rect 981 1503 983 1507
rect 968 1502 973 1503
rect 978 1502 983 1503
rect 456 1403 458 1407
rect 458 1403 461 1407
rect 466 1403 469 1407
rect 469 1403 471 1407
rect 456 1402 461 1403
rect 466 1402 471 1403
rect 1480 1403 1482 1407
rect 1482 1403 1485 1407
rect 1490 1403 1493 1407
rect 1493 1403 1495 1407
rect 1480 1402 1485 1403
rect 1490 1402 1495 1403
rect 968 1303 970 1307
rect 970 1303 973 1307
rect 978 1303 981 1307
rect 981 1303 983 1307
rect 968 1302 973 1303
rect 978 1302 983 1303
rect 456 1203 458 1207
rect 458 1203 461 1207
rect 466 1203 469 1207
rect 469 1203 471 1207
rect 456 1202 461 1203
rect 466 1202 471 1203
rect 1480 1203 1482 1207
rect 1482 1203 1485 1207
rect 1490 1203 1493 1207
rect 1493 1203 1495 1207
rect 1480 1202 1485 1203
rect 1490 1202 1495 1203
rect 968 1103 970 1107
rect 970 1103 973 1107
rect 978 1103 981 1107
rect 981 1103 983 1107
rect 968 1102 973 1103
rect 978 1102 983 1103
rect 456 1003 458 1007
rect 458 1003 461 1007
rect 466 1003 469 1007
rect 469 1003 471 1007
rect 456 1002 461 1003
rect 466 1002 471 1003
rect 1480 1003 1482 1007
rect 1482 1003 1485 1007
rect 1490 1003 1493 1007
rect 1493 1003 1495 1007
rect 1480 1002 1485 1003
rect 1490 1002 1495 1003
rect 968 903 970 907
rect 970 903 973 907
rect 978 903 981 907
rect 981 903 983 907
rect 968 902 973 903
rect 978 902 983 903
rect 456 803 458 807
rect 458 803 461 807
rect 466 803 469 807
rect 469 803 471 807
rect 456 802 461 803
rect 466 802 471 803
rect 1480 803 1482 807
rect 1482 803 1485 807
rect 1490 803 1493 807
rect 1493 803 1495 807
rect 1480 802 1485 803
rect 1490 802 1495 803
rect 968 703 970 707
rect 970 703 973 707
rect 978 703 981 707
rect 981 703 983 707
rect 968 702 973 703
rect 978 702 983 703
rect 456 603 458 607
rect 458 603 461 607
rect 466 603 469 607
rect 469 603 471 607
rect 456 602 461 603
rect 466 602 471 603
rect 1480 603 1482 607
rect 1482 603 1485 607
rect 1490 603 1493 607
rect 1493 603 1495 607
rect 1480 602 1485 603
rect 1490 602 1495 603
rect 968 503 970 507
rect 970 503 973 507
rect 978 503 981 507
rect 981 503 983 507
rect 968 502 973 503
rect 978 502 983 503
rect 456 403 458 407
rect 458 403 461 407
rect 466 403 469 407
rect 469 403 471 407
rect 456 402 461 403
rect 466 402 471 403
rect 1480 403 1482 407
rect 1482 403 1485 407
rect 1490 403 1493 407
rect 1493 403 1495 407
rect 1480 402 1485 403
rect 1490 402 1495 403
rect 968 303 970 307
rect 970 303 973 307
rect 978 303 981 307
rect 981 303 983 307
rect 968 302 973 303
rect 978 302 983 303
rect 456 203 458 207
rect 458 203 461 207
rect 466 203 469 207
rect 469 203 471 207
rect 456 202 461 203
rect 466 202 471 203
rect 1480 203 1482 207
rect 1482 203 1485 207
rect 1490 203 1493 207
rect 1493 203 1495 207
rect 1480 202 1485 203
rect 1490 202 1495 203
rect 968 103 970 107
rect 970 103 973 107
rect 978 103 981 107
rect 981 103 983 107
rect 968 102 973 103
rect 978 102 983 103
rect 456 3 458 7
rect 458 3 461 7
rect 466 3 469 7
rect 469 3 471 7
rect 456 2 461 3
rect 466 2 471 3
rect 1480 3 1482 7
rect 1482 3 1485 7
rect 1490 3 1493 7
rect 1493 3 1495 7
rect 1480 2 1485 3
rect 1490 2 1495 3
<< metal6 >>
rect 456 1607 472 1730
rect 461 1602 466 1607
rect 471 1602 472 1607
rect 456 1407 472 1602
rect 461 1402 466 1407
rect 471 1402 472 1407
rect 456 1207 472 1402
rect 461 1202 466 1207
rect 471 1202 472 1207
rect 456 1007 472 1202
rect 461 1002 466 1007
rect 471 1002 472 1007
rect 456 807 472 1002
rect 461 802 466 807
rect 471 802 472 807
rect 456 607 472 802
rect 461 602 466 607
rect 471 602 472 607
rect 456 407 472 602
rect 461 402 466 407
rect 471 402 472 407
rect 456 207 472 402
rect 461 202 466 207
rect 471 202 472 207
rect 456 7 472 202
rect 461 2 466 7
rect 471 2 472 7
rect 456 -30 472 2
rect 968 1707 984 1730
rect 973 1702 978 1707
rect 983 1702 984 1707
rect 968 1507 984 1702
rect 973 1502 978 1507
rect 983 1502 984 1507
rect 968 1307 984 1502
rect 973 1302 978 1307
rect 983 1302 984 1307
rect 968 1107 984 1302
rect 973 1102 978 1107
rect 983 1102 984 1107
rect 968 907 984 1102
rect 973 902 978 907
rect 983 902 984 907
rect 968 707 984 902
rect 973 702 978 707
rect 983 702 984 707
rect 968 507 984 702
rect 973 502 978 507
rect 983 502 984 507
rect 968 307 984 502
rect 973 302 978 307
rect 983 302 984 307
rect 968 107 984 302
rect 973 102 978 107
rect 983 102 984 107
rect 968 -30 984 102
rect 1480 1607 1496 1730
rect 1485 1602 1490 1607
rect 1495 1602 1496 1607
rect 1480 1407 1496 1602
rect 1485 1402 1490 1407
rect 1495 1402 1496 1407
rect 1480 1207 1496 1402
rect 1485 1202 1490 1207
rect 1495 1202 1496 1207
rect 1480 1007 1496 1202
rect 1485 1002 1490 1007
rect 1495 1002 1496 1007
rect 1480 807 1496 1002
rect 1485 802 1490 807
rect 1495 802 1496 807
rect 1480 607 1496 802
rect 1485 602 1490 607
rect 1495 602 1496 607
rect 1480 407 1496 602
rect 1485 402 1490 407
rect 1495 402 1496 407
rect 1480 207 1496 402
rect 1485 202 1490 207
rect 1495 202 1496 207
rect 1480 7 1496 202
rect 1485 2 1490 7
rect 1495 2 1496 7
rect 1480 -30 1496 2
use INVX1  INVX1_6
timestamp 1696677024
transform 1 0 4 0 -1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_8
timestamp 1696677024
transform 1 0 20 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_9
timestamp 1696677024
transform -1 0 76 0 -1 105
box -2 -3 26 103
use NOR3X1  NOR3X1_1
timestamp 1696677024
transform -1 0 140 0 -1 105
box -2 -3 66 103
use BUFX2  BUFX2_17
timestamp 1696677024
transform -1 0 28 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_14
timestamp 1696677024
transform -1 0 124 0 1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_6
timestamp 1696677024
transform -1 0 164 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_2
timestamp 1696677024
transform -1 0 188 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_9
timestamp 1696677024
transform -1 0 220 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_8
timestamp 1696677024
transform -1 0 148 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_29
timestamp 1696677024
transform 1 0 148 0 1 105
box -2 -3 98 103
use INVX2  INVX2_16
timestamp 1696677024
transform 1 0 220 0 -1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_7
timestamp 1696677024
transform 1 0 236 0 -1 105
box -2 -3 26 103
use NOR3X1  NOR3X1_2
timestamp 1696677024
transform -1 0 324 0 -1 105
box -2 -3 66 103
use NOR2X1  NOR2X1_10
timestamp 1696677024
transform -1 0 268 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_8
timestamp 1696677024
transform 1 0 268 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_58
timestamp 1696677024
transform 1 0 300 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_59
timestamp 1696677024
transform -1 0 348 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_16
timestamp 1696677024
transform -1 0 444 0 -1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_106
timestamp 1696677024
transform 1 0 324 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_30
timestamp 1696677024
transform -1 0 444 0 1 105
box -2 -3 98 103
use FILL  FILL_0_0_0
timestamp 1696677024
transform 1 0 444 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_0_1
timestamp 1696677024
transform 1 0 452 0 -1 105
box -2 -3 10 103
use OAI21X1  OAI21X1_10
timestamp 1696677024
transform 1 0 460 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_11
timestamp 1696677024
transform 1 0 492 0 -1 105
box -2 -3 26 103
use FILL  FILL_1_0_0
timestamp 1696677024
transform 1 0 444 0 1 105
box -2 -3 10 103
use FILL  FILL_1_0_1
timestamp 1696677024
transform 1 0 452 0 1 105
box -2 -3 10 103
use AND2X2  AND2X2_2
timestamp 1696677024
transform 1 0 460 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_31
timestamp 1696677024
transform -1 0 588 0 1 105
box -2 -3 98 103
use INVX1  INVX1_5
timestamp 1696677024
transform 1 0 516 0 -1 105
box -2 -3 18 103
use OAI21X1  OAI21X1_7
timestamp 1696677024
transform 1 0 532 0 -1 105
box -2 -3 34 103
use BUFX2  BUFX2_32
timestamp 1696677024
transform 1 0 564 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_7
timestamp 1696677024
transform 1 0 588 0 -1 105
box -2 -3 34 103
use CLKBUF1  CLKBUF1_7
timestamp 1696677024
transform -1 0 660 0 1 105
box -2 -3 74 103
use NAND2X1  NAND2X1_60
timestamp 1696677024
transform 1 0 620 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_11
timestamp 1696677024
transform 1 0 644 0 -1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_26
timestamp 1696677024
transform 1 0 660 0 1 105
box -2 -3 98 103
use INVX1  INVX1_2
timestamp 1696677024
transform 1 0 740 0 -1 105
box -2 -3 18 103
use AOI21X1  AOI21X1_5
timestamp 1696677024
transform 1 0 756 0 -1 105
box -2 -3 34 103
use OR2X2  OR2X2_1
timestamp 1696677024
transform 1 0 788 0 -1 105
box -2 -3 34 103
use AND2X2  AND2X2_1
timestamp 1696677024
transform -1 0 788 0 1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_57
timestamp 1696677024
transform -1 0 812 0 1 105
box -2 -3 26 103
use INVX1  INVX1_4
timestamp 1696677024
transform 1 0 820 0 -1 105
box -2 -3 18 103
use NAND3X1  NAND3X1_1
timestamp 1696677024
transform 1 0 836 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_54
timestamp 1696677024
transform -1 0 892 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_22
timestamp 1696677024
transform 1 0 892 0 -1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_107
timestamp 1696677024
transform -1 0 836 0 1 105
box -2 -3 26 103
use INVX1  INVX1_3
timestamp 1696677024
transform 1 0 836 0 1 105
box -2 -3 18 103
use AOI21X1  AOI21X1_6
timestamp 1696677024
transform 1 0 852 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_6
timestamp 1696677024
transform -1 0 916 0 1 105
box -2 -3 34 103
use FILL  FILL_0_1_0
timestamp 1696677024
transform 1 0 988 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_1_1
timestamp 1696677024
transform 1 0 996 0 -1 105
box -2 -3 10 103
use NOR2X1  NOR2X1_102
timestamp 1696677024
transform 1 0 1004 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_105
timestamp 1696677024
transform -1 0 940 0 1 105
box -2 -3 26 103
use BUFX2  BUFX2_49
timestamp 1696677024
transform 1 0 940 0 1 105
box -2 -3 26 103
use FILL  FILL_1_1_0
timestamp 1696677024
transform 1 0 964 0 1 105
box -2 -3 10 103
use FILL  FILL_1_1_1
timestamp 1696677024
transform 1 0 972 0 1 105
box -2 -3 10 103
use NOR3X1  NOR3X1_13
timestamp 1696677024
transform 1 0 980 0 1 105
box -2 -3 66 103
use NAND2X1  NAND2X1_50
timestamp 1696677024
transform -1 0 1052 0 -1 105
box -2 -3 26 103
use AND2X2  AND2X2_19
timestamp 1696677024
transform -1 0 1084 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_7
timestamp 1696677024
transform -1 0 1180 0 -1 105
box -2 -3 98 103
use NAND2X1  NAND2X1_56
timestamp 1696677024
transform 1 0 1044 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_5
timestamp 1696677024
transform 1 0 1068 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_5
timestamp 1696677024
transform 1 0 1100 0 1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_1
timestamp 1696677024
transform -1 0 1204 0 -1 105
box -2 -3 26 103
use NOR2X1  NOR2X1_2
timestamp 1696677024
transform -1 0 1228 0 -1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_4
timestamp 1696677024
transform -1 0 1156 0 1 105
box -2 -3 34 103
use INVX2  INVX2_1
timestamp 1696677024
transform -1 0 1172 0 1 105
box -2 -3 18 103
use NOR2X1  NOR2X1_3
timestamp 1696677024
transform -1 0 1196 0 1 105
box -2 -3 26 103
use INVX1  INVX1_1
timestamp 1696677024
transform -1 0 1212 0 1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_23
timestamp 1696677024
transform -1 0 1308 0 1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_2
timestamp 1696677024
transform 1 0 1228 0 -1 105
box -2 -3 34 103
use NAND2X1  NAND2X1_51
timestamp 1696677024
transform 1 0 1260 0 -1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_8
timestamp 1696677024
transform 1 0 1284 0 -1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_4
timestamp 1696677024
transform 1 0 1308 0 1 105
box -2 -3 26 103
use AND2X2  AND2X2_20
timestamp 1696677024
transform 1 0 1380 0 -1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_24
timestamp 1696677024
transform 1 0 1412 0 -1 105
box -2 -3 98 103
use OAI21X1  OAI21X1_3
timestamp 1696677024
transform -1 0 1364 0 1 105
box -2 -3 34 103
use OAI21X1  OAI21X1_4
timestamp 1696677024
transform 1 0 1364 0 1 105
box -2 -3 34 103
use AOI21X1  AOI21X1_3
timestamp 1696677024
transform 1 0 1396 0 1 105
box -2 -3 34 103
use FILL  FILL_0_2_0
timestamp 1696677024
transform -1 0 1516 0 -1 105
box -2 -3 10 103
use FILL  FILL_0_2_1
timestamp 1696677024
transform -1 0 1524 0 -1 105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_17
timestamp 1696677024
transform 1 0 1428 0 1 105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_9
timestamp 1696677024
transform -1 0 1620 0 -1 105
box -2 -3 98 103
use FILL  FILL_1_2_0
timestamp 1696677024
transform 1 0 1524 0 1 105
box -2 -3 10 103
use FILL  FILL_1_2_1
timestamp 1696677024
transform 1 0 1532 0 1 105
box -2 -3 10 103
use INVX2  INVX2_15
timestamp 1696677024
transform 1 0 1540 0 1 105
box -2 -3 18 103
use OR2X2  OR2X2_10
timestamp 1696677024
transform -1 0 1588 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_21
timestamp 1696677024
transform 1 0 1588 0 1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_103
timestamp 1696677024
transform 1 0 1620 0 -1 105
box -2 -3 26 103
use BUFX2  BUFX2_41
timestamp 1696677024
transform 1 0 1644 0 -1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_1
timestamp 1696677024
transform 1 0 1668 0 -1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_1
timestamp 1696677024
transform 1 0 1700 0 -1 105
box -2 -3 26 103
use NAND2X1  NAND2X1_53
timestamp 1696677024
transform -1 0 1708 0 1 105
box -2 -3 26 103
use AOI21X1  AOI21X1_2
timestamp 1696677024
transform -1 0 1740 0 1 105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_6
timestamp 1696677024
transform -1 0 1820 0 -1 105
box -2 -3 98 103
use NOR2X1  NOR2X1_57
timestamp 1696677024
transform -1 0 1844 0 -1 105
box -2 -3 26 103
use INVX2  INVX2_17
timestamp 1696677024
transform -1 0 1756 0 1 105
box -2 -3 18 103
use NAND2X1  NAND2X1_52
timestamp 1696677024
transform -1 0 1780 0 1 105
box -2 -3 26 103
use OAI21X1  OAI21X1_67
timestamp 1696677024
transform -1 0 1812 0 1 105
box -2 -3 34 103
use NOR2X1  NOR2X1_108
timestamp 1696677024
transform -1 0 1836 0 1 105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_3
timestamp 1696677024
transform 1 0 1844 0 -1 105
box -2 -3 98 103
use INVX1  INVX1_23
timestamp 1696677024
transform 1 0 1836 0 1 105
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_18
timestamp 1696677024
transform 1 0 1852 0 1 105
box -2 -3 98 103
use FILL  FILL_1_1
timestamp 1696677024
transform -1 0 1948 0 -1 105
box -2 -3 10 103
use FILL  FILL_1_2
timestamp 1696677024
transform -1 0 1956 0 -1 105
box -2 -3 10 103
use FILL  FILL_2_1
timestamp 1696677024
transform 1 0 1948 0 1 105
box -2 -3 10 103
use OR2X2  OR2X2_5
timestamp 1696677024
transform 1 0 4 0 -1 305
box -2 -3 34 103
use OR2X2  OR2X2_4
timestamp 1696677024
transform 1 0 36 0 -1 305
box -2 -3 34 103
use INVX1  INVX1_31
timestamp 1696677024
transform 1 0 68 0 -1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_13
timestamp 1696677024
transform 1 0 84 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_28
timestamp 1696677024
transform 1 0 180 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_15
timestamp 1696677024
transform 1 0 276 0 -1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_98
timestamp 1696677024
transform -1 0 396 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_77
timestamp 1696677024
transform 1 0 396 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_0_0
timestamp 1696677024
transform 1 0 492 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_0_1
timestamp 1696677024
transform 1 0 500 0 -1 305
box -2 -3 10 103
use AND2X2  AND2X2_5
timestamp 1696677024
transform 1 0 508 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_96
timestamp 1696677024
transform -1 0 636 0 -1 305
box -2 -3 98 103
use BUFX2  BUFX2_54
timestamp 1696677024
transform -1 0 660 0 -1 305
box -2 -3 26 103
use OR2X2  OR2X2_8
timestamp 1696677024
transform -1 0 692 0 -1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_68
timestamp 1696677024
transform 1 0 692 0 -1 305
box -2 -3 26 103
use INVX1  INVX1_34
timestamp 1696677024
transform 1 0 716 0 -1 305
box -2 -3 18 103
use NAND3X1  NAND3X1_22
timestamp 1696677024
transform 1 0 732 0 -1 305
box -2 -3 34 103
use INVX2  INVX2_14
timestamp 1696677024
transform 1 0 764 0 -1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_12
timestamp 1696677024
transform -1 0 876 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_27
timestamp 1696677024
transform -1 0 972 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_1_0
timestamp 1696677024
transform 1 0 972 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_1_1
timestamp 1696677024
transform 1 0 980 0 -1 305
box -2 -3 10 103
use AND2X2  AND2X2_6
timestamp 1696677024
transform 1 0 988 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_25
timestamp 1696677024
transform -1 0 1116 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_10
timestamp 1696677024
transform -1 0 1212 0 -1 305
box -2 -3 98 103
use INVX1  INVX1_29
timestamp 1696677024
transform 1 0 1212 0 -1 305
box -2 -3 18 103
use CLKBUF1  CLKBUF1_6
timestamp 1696677024
transform -1 0 1300 0 -1 305
box -2 -3 74 103
use INVX1  INVX1_30
timestamp 1696677024
transform 1 0 1300 0 -1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_65
timestamp 1696677024
transform 1 0 1316 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_32
timestamp 1696677024
transform 1 0 1340 0 -1 305
box -2 -3 98 103
use FILL  FILL_2_2_0
timestamp 1696677024
transform 1 0 1436 0 -1 305
box -2 -3 10 103
use FILL  FILL_2_2_1
timestamp 1696677024
transform 1 0 1444 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_2
timestamp 1696677024
transform 1 0 1452 0 -1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_1
timestamp 1696677024
transform 1 0 1548 0 -1 305
box -2 -3 98 103
use OAI21X1  OAI21X1_68
timestamp 1696677024
transform -1 0 1676 0 -1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_5
timestamp 1696677024
transform -1 0 1772 0 -1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_109
timestamp 1696677024
transform 1 0 1772 0 -1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_4
timestamp 1696677024
transform 1 0 1796 0 -1 305
box -2 -3 98 103
use BUFX2  BUFX2_48
timestamp 1696677024
transform -1 0 1916 0 -1 305
box -2 -3 26 103
use BUFX2  BUFX2_34
timestamp 1696677024
transform 1 0 1916 0 -1 305
box -2 -3 26 103
use FILL  FILL_3_1
timestamp 1696677024
transform -1 0 1948 0 -1 305
box -2 -3 10 103
use FILL  FILL_3_2
timestamp 1696677024
transform -1 0 1956 0 -1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_46
timestamp 1696677024
transform -1 0 100 0 1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_62
timestamp 1696677024
transform -1 0 196 0 1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_49
timestamp 1696677024
transform 1 0 196 0 1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_93
timestamp 1696677024
transform -1 0 388 0 1 305
box -2 -3 98 103
use AND2X2  AND2X2_17
timestamp 1696677024
transform 1 0 388 0 1 305
box -2 -3 34 103
use OAI22X1  OAI22X1_4
timestamp 1696677024
transform 1 0 420 0 1 305
box -2 -3 42 103
use FILL  FILL_3_0_0
timestamp 1696677024
transform -1 0 468 0 1 305
box -2 -3 10 103
use FILL  FILL_3_0_1
timestamp 1696677024
transform -1 0 476 0 1 305
box -2 -3 10 103
use AND2X2  AND2X2_18
timestamp 1696677024
transform -1 0 508 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_99
timestamp 1696677024
transform -1 0 532 0 1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_80
timestamp 1696677024
transform -1 0 628 0 1 305
box -2 -3 98 103
use OR2X2  OR2X2_6
timestamp 1696677024
transform -1 0 660 0 1 305
box -2 -3 34 103
use INVX1  INVX1_32
timestamp 1696677024
transform 1 0 660 0 1 305
box -2 -3 18 103
use NOR2X1  NOR2X1_66
timestamp 1696677024
transform 1 0 676 0 1 305
box -2 -3 26 103
use NAND2X1  NAND2X1_31
timestamp 1696677024
transform -1 0 724 0 1 305
box -2 -3 26 103
use AND2X2  AND2X2_7
timestamp 1696677024
transform -1 0 756 0 1 305
box -2 -3 34 103
use NOR2X1  NOR2X1_67
timestamp 1696677024
transform 1 0 756 0 1 305
box -2 -3 26 103
use INVX1  INVX1_19
timestamp 1696677024
transform 1 0 780 0 1 305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_115
timestamp 1696677024
transform 1 0 796 0 1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_118
timestamp 1696677024
transform 1 0 892 0 1 305
box -2 -3 98 103
use FILL  FILL_3_1_0
timestamp 1696677024
transform -1 0 996 0 1 305
box -2 -3 10 103
use FILL  FILL_3_1_1
timestamp 1696677024
transform -1 0 1004 0 1 305
box -2 -3 10 103
use AND2X2  AND2X2_9
timestamp 1696677024
transform -1 0 1036 0 1 305
box -2 -3 34 103
use NOR3X1  NOR3X1_7
timestamp 1696677024
transform 1 0 1036 0 1 305
box -2 -3 66 103
use NOR2X1  NOR2X1_104
timestamp 1696677024
transform -1 0 1124 0 1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_117
timestamp 1696677024
transform -1 0 1220 0 1 305
box -2 -3 98 103
use NOR2X1  NOR2X1_64
timestamp 1696677024
transform 1 0 1220 0 1 305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_116
timestamp 1696677024
transform -1 0 1340 0 1 305
box -2 -3 98 103
use BUFX2  BUFX2_38
timestamp 1696677024
transform -1 0 1364 0 1 305
box -2 -3 26 103
use BUFX2  BUFX2_39
timestamp 1696677024
transform 1 0 1364 0 1 305
box -2 -3 26 103
use CLKBUF1  CLKBUF1_4
timestamp 1696677024
transform 1 0 1388 0 1 305
box -2 -3 74 103
use FILL  FILL_3_2_0
timestamp 1696677024
transform 1 0 1460 0 1 305
box -2 -3 10 103
use FILL  FILL_3_2_1
timestamp 1696677024
transform 1 0 1468 0 1 305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_106
timestamp 1696677024
transform 1 0 1476 0 1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_110
timestamp 1696677024
transform 1 0 1572 0 1 305
box -2 -3 98 103
use AOI21X1  AOI21X1_1
timestamp 1696677024
transform -1 0 1700 0 1 305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_20
timestamp 1696677024
transform -1 0 1796 0 1 305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_19
timestamp 1696677024
transform 1 0 1796 0 1 305
box -2 -3 98 103
use BUFX2  BUFX2_47
timestamp 1696677024
transform 1 0 1892 0 1 305
box -2 -3 26 103
use BUFX2  BUFX2_36
timestamp 1696677024
transform 1 0 1916 0 1 305
box -2 -3 26 103
use FILL  FILL_4_1
timestamp 1696677024
transform 1 0 1940 0 1 305
box -2 -3 10 103
use FILL  FILL_4_2
timestamp 1696677024
transform 1 0 1948 0 1 305
box -2 -3 10 103
use BUFX2  BUFX2_25
timestamp 1696677024
transform -1 0 28 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_33
timestamp 1696677024
transform -1 0 124 0 -1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_17
timestamp 1696677024
transform -1 0 148 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_35
timestamp 1696677024
transform 1 0 148 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_51
timestamp 1696677024
transform 1 0 244 0 -1 505
box -2 -3 98 103
use NOR3X1  NOR3X1_12
timestamp 1696677024
transform -1 0 404 0 -1 505
box -2 -3 66 103
use XOR2X1  XOR2X1_7
timestamp 1696677024
transform -1 0 460 0 -1 505
box -2 -3 58 103
use FILL  FILL_4_0_0
timestamp 1696677024
transform -1 0 468 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_0_1
timestamp 1696677024
transform -1 0 476 0 -1 505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_50
timestamp 1696677024
transform -1 0 572 0 -1 505
box -2 -3 98 103
use CLKBUF1  CLKBUF1_8
timestamp 1696677024
transform -1 0 644 0 -1 505
box -2 -3 74 103
use BUFX2  BUFX2_52
timestamp 1696677024
transform -1 0 668 0 -1 505
box -2 -3 26 103
use INVX1  INVX1_27
timestamp 1696677024
transform -1 0 684 0 -1 505
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_34
timestamp 1696677024
transform -1 0 780 0 -1 505
box -2 -3 98 103
use OAI21X1  OAI21X1_39
timestamp 1696677024
transform -1 0 812 0 -1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_23
timestamp 1696677024
transform 1 0 812 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_48
timestamp 1696677024
transform -1 0 860 0 -1 505
box -2 -3 26 103
use INVX2  INVX2_9
timestamp 1696677024
transform -1 0 876 0 -1 505
box -2 -3 18 103
use NOR2X1  NOR2X1_45
timestamp 1696677024
transform 1 0 876 0 -1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_21
timestamp 1696677024
transform 1 0 900 0 -1 505
box -2 -3 26 103
use INVX2  INVX2_8
timestamp 1696677024
transform 1 0 924 0 -1 505
box -2 -3 18 103
use FILL  FILL_4_1_0
timestamp 1696677024
transform -1 0 948 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_1_1
timestamp 1696677024
transform -1 0 956 0 -1 505
box -2 -3 10 103
use NOR3X1  NOR3X1_8
timestamp 1696677024
transform -1 0 1020 0 -1 505
box -2 -3 66 103
use INVX1  INVX1_33
timestamp 1696677024
transform -1 0 1036 0 -1 505
box -2 -3 18 103
use BUFX2  BUFX2_53
timestamp 1696677024
transform 1 0 1036 0 -1 505
box -2 -3 26 103
use NOR3X1  NOR3X1_6
timestamp 1696677024
transform 1 0 1060 0 -1 505
box -2 -3 66 103
use AOI22X1  AOI22X1_1
timestamp 1696677024
transform 1 0 1124 0 -1 505
box -2 -3 42 103
use AOI21X1  AOI21X1_30
timestamp 1696677024
transform 1 0 1164 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_113
timestamp 1696677024
transform -1 0 1292 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_107
timestamp 1696677024
transform 1 0 1292 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_111
timestamp 1696677024
transform -1 0 1484 0 -1 505
box -2 -3 98 103
use FILL  FILL_4_2_0
timestamp 1696677024
transform 1 0 1484 0 -1 505
box -2 -3 10 103
use FILL  FILL_4_2_1
timestamp 1696677024
transform 1 0 1492 0 -1 505
box -2 -3 10 103
use NOR2X1  NOR2X1_62
timestamp 1696677024
transform 1 0 1500 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_61
timestamp 1696677024
transform 1 0 1524 0 -1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_20
timestamp 1696677024
transform -1 0 1580 0 -1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_105
timestamp 1696677024
transform -1 0 1676 0 -1 505
box -2 -3 98 103
use NAND2X1  NAND2X1_27
timestamp 1696677024
transform -1 0 1700 0 -1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_59
timestamp 1696677024
transform 1 0 1700 0 -1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_109
timestamp 1696677024
transform 1 0 1724 0 -1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_101
timestamp 1696677024
transform 1 0 1820 0 -1 505
box -2 -3 98 103
use BUFX2  BUFX2_44
timestamp 1696677024
transform 1 0 1916 0 -1 505
box -2 -3 26 103
use FILL  FILL_5_1
timestamp 1696677024
transform -1 0 1948 0 -1 505
box -2 -3 10 103
use FILL  FILL_5_2
timestamp 1696677024
transform -1 0 1956 0 -1 505
box -2 -3 10 103
use CLKBUF1  CLKBUF1_13
timestamp 1696677024
transform 1 0 4 0 1 505
box -2 -3 74 103
use NOR2X1  NOR2X1_20
timestamp 1696677024
transform 1 0 76 0 1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_9
timestamp 1696677024
transform 1 0 100 0 1 505
box -2 -3 50 103
use NAND2X1  NAND2X1_46
timestamp 1696677024
transform 1 0 148 0 1 505
box -2 -3 26 103
use BUFX4  BUFX4_7
timestamp 1696677024
transform -1 0 204 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_22
timestamp 1696677024
transform 1 0 204 0 1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_11
timestamp 1696677024
transform 1 0 228 0 1 505
box -2 -3 50 103
use NAND2X1  NAND2X1_48
timestamp 1696677024
transform 1 0 276 0 1 505
box -2 -3 26 103
use XOR2X1  XOR2X1_8
timestamp 1696677024
transform 1 0 300 0 1 505
box -2 -3 58 103
use INVX1  INVX1_54
timestamp 1696677024
transform 1 0 356 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_62
timestamp 1696677024
transform 1 0 372 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_47
timestamp 1696677024
transform -1 0 428 0 1 505
box -2 -3 26 103
use INVX1  INVX1_56
timestamp 1696677024
transform 1 0 428 0 1 505
box -2 -3 18 103
use FILL  FILL_5_0_0
timestamp 1696677024
transform 1 0 444 0 1 505
box -2 -3 10 103
use FILL  FILL_5_0_1
timestamp 1696677024
transform 1 0 452 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_64
timestamp 1696677024
transform 1 0 460 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_49
timestamp 1696677024
transform 1 0 492 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_36
timestamp 1696677024
transform -1 0 612 0 1 505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_52
timestamp 1696677024
transform -1 0 708 0 1 505
box -2 -3 98 103
use NOR2X1  NOR2X1_23
timestamp 1696677024
transform 1 0 708 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_21
timestamp 1696677024
transform 1 0 732 0 1 505
box -2 -3 26 103
use MUX2X1  MUX2X1_12
timestamp 1696677024
transform 1 0 756 0 1 505
box -2 -3 50 103
use AOI22X1  AOI22X1_3
timestamp 1696677024
transform 1 0 804 0 1 505
box -2 -3 42 103
use AOI21X1  AOI21X1_32
timestamp 1696677024
transform -1 0 876 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_47
timestamp 1696677024
transform 1 0 876 0 1 505
box -2 -3 26 103
use NAND2X1  NAND2X1_22
timestamp 1696677024
transform 1 0 900 0 1 505
box -2 -3 26 103
use INVX1  INVX1_18
timestamp 1696677024
transform 1 0 924 0 1 505
box -2 -3 18 103
use FILL  FILL_5_1_0
timestamp 1696677024
transform 1 0 940 0 1 505
box -2 -3 10 103
use FILL  FILL_5_1_1
timestamp 1696677024
transform 1 0 948 0 1 505
box -2 -3 10 103
use NOR3X1  NOR3X1_5
timestamp 1696677024
transform 1 0 956 0 1 505
box -2 -3 66 103
use AOI22X1  AOI22X1_4
timestamp 1696677024
transform 1 0 1020 0 1 505
box -2 -3 42 103
use NOR2X1  NOR2X1_46
timestamp 1696677024
transform -1 0 1084 0 1 505
box -2 -3 26 103
use AND2X2  AND2X2_4
timestamp 1696677024
transform 1 0 1084 0 1 505
box -2 -3 34 103
use AOI22X1  AOI22X1_2
timestamp 1696677024
transform -1 0 1156 0 1 505
box -2 -3 42 103
use OR2X2  OR2X2_9
timestamp 1696677024
transform -1 0 1188 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_31
timestamp 1696677024
transform 1 0 1188 0 1 505
box -2 -3 34 103
use BUFX2  BUFX2_55
timestamp 1696677024
transform 1 0 1220 0 1 505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_114
timestamp 1696677024
transform -1 0 1340 0 1 505
box -2 -3 98 103
use AOI21X1  AOI21X1_29
timestamp 1696677024
transform -1 0 1372 0 1 505
box -2 -3 34 103
use AOI21X1  AOI21X1_28
timestamp 1696677024
transform -1 0 1404 0 1 505
box -2 -3 34 103
use INVX1  INVX1_25
timestamp 1696677024
transform 1 0 1404 0 1 505
box -2 -3 18 103
use NAND2X1  NAND2X1_29
timestamp 1696677024
transform 1 0 1420 0 1 505
box -2 -3 26 103
use AOI21X1  AOI21X1_27
timestamp 1696677024
transform 1 0 1444 0 1 505
box -2 -3 34 103
use FILL  FILL_5_2_0
timestamp 1696677024
transform -1 0 1484 0 1 505
box -2 -3 10 103
use FILL  FILL_5_2_1
timestamp 1696677024
transform -1 0 1492 0 1 505
box -2 -3 10 103
use OAI21X1  OAI21X1_45
timestamp 1696677024
transform -1 0 1524 0 1 505
box -2 -3 34 103
use INVX2  INVX2_13
timestamp 1696677024
transform 1 0 1524 0 1 505
box -2 -3 18 103
use XNOR2X1  XNOR2X1_7
timestamp 1696677024
transform -1 0 1596 0 1 505
box -2 -3 58 103
use NOR2X1  NOR2X1_56
timestamp 1696677024
transform -1 0 1620 0 1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_19
timestamp 1696677024
transform -1 0 1652 0 1 505
box -2 -3 34 103
use NAND2X1  NAND2X1_28
timestamp 1696677024
transform 1 0 1652 0 1 505
box -2 -3 26 103
use NOR2X1  NOR2X1_60
timestamp 1696677024
transform 1 0 1676 0 1 505
box -2 -3 26 103
use NAND3X1  NAND3X1_21
timestamp 1696677024
transform 1 0 1700 0 1 505
box -2 -3 34 103
use INVX1  INVX1_24
timestamp 1696677024
transform 1 0 1732 0 1 505
box -2 -3 18 103
use OAI21X1  OAI21X1_44
timestamp 1696677024
transform -1 0 1780 0 1 505
box -2 -3 34 103
use NOR2X1  NOR2X1_58
timestamp 1696677024
transform 1 0 1780 0 1 505
box -2 -3 26 103
use OAI21X1  OAI21X1_43
timestamp 1696677024
transform -1 0 1836 0 1 505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_97
timestamp 1696677024
transform 1 0 1836 0 1 505
box -2 -3 98 103
use INVX1  INVX1_45
timestamp 1696677024
transform -1 0 1948 0 1 505
box -2 -3 18 103
use FILL  FILL_6_1
timestamp 1696677024
transform 1 0 1948 0 1 505
box -2 -3 10 103
use BUFX2  BUFX2_24
timestamp 1696677024
transform -1 0 28 0 -1 705
box -2 -3 26 103
use CLKBUF1  CLKBUF1_9
timestamp 1696677024
transform 1 0 28 0 -1 705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_64
timestamp 1696677024
transform -1 0 196 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_61
timestamp 1696677024
transform -1 0 228 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_53
timestamp 1696677024
transform -1 0 244 0 -1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_54
timestamp 1696677024
transform 1 0 244 0 -1 705
box -2 -3 98 103
use OAI21X1  OAI21X1_63
timestamp 1696677024
transform -1 0 372 0 -1 705
box -2 -3 34 103
use INVX1  INVX1_55
timestamp 1696677024
transform -1 0 388 0 -1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_78
timestamp 1696677024
transform 1 0 388 0 -1 705
box -2 -3 98 103
use FILL  FILL_6_0_0
timestamp 1696677024
transform 1 0 484 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_0_1
timestamp 1696677024
transform 1 0 492 0 -1 705
box -2 -3 10 103
use INVX1  INVX1_9
timestamp 1696677024
transform 1 0 500 0 -1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_8
timestamp 1696677024
transform -1 0 540 0 -1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_12
timestamp 1696677024
transform 1 0 540 0 -1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_16
timestamp 1696677024
transform -1 0 604 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_33
timestamp 1696677024
transform -1 0 628 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_79
timestamp 1696677024
transform -1 0 724 0 -1 705
box -2 -3 98 103
use MUX2X1  MUX2X1_10
timestamp 1696677024
transform 1 0 724 0 -1 705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_138
timestamp 1696677024
transform -1 0 868 0 -1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_80
timestamp 1696677024
transform 1 0 868 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_122
timestamp 1696677024
transform 1 0 892 0 -1 705
box -2 -3 98 103
use FILL  FILL_6_1_0
timestamp 1696677024
transform -1 0 996 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_1_1
timestamp 1696677024
transform -1 0 1004 0 -1 705
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_131
timestamp 1696677024
transform -1 0 1100 0 -1 705
box -2 -3 98 103
use INVX1  INVX1_28
timestamp 1696677024
transform 1 0 1100 0 -1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_63
timestamp 1696677024
transform 1 0 1116 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_149
timestamp 1696677024
transform 1 0 1140 0 -1 705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_12
timestamp 1696677024
transform 1 0 1236 0 -1 705
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_112
timestamp 1696677024
transform 1 0 1308 0 -1 705
box -2 -3 98 103
use CLKBUF1  CLKBUF1_14
timestamp 1696677024
transform 1 0 1404 0 -1 705
box -2 -3 74 103
use FILL  FILL_6_2_0
timestamp 1696677024
transform -1 0 1484 0 -1 705
box -2 -3 10 103
use FILL  FILL_6_2_1
timestamp 1696677024
transform -1 0 1492 0 -1 705
box -2 -3 10 103
use BUFX2  BUFX2_50
timestamp 1696677024
transform -1 0 1516 0 -1 705
box -2 -3 26 103
use AND2X2  AND2X2_8
timestamp 1696677024
transform -1 0 1548 0 -1 705
box -2 -3 34 103
use BUFX2  BUFX2_56
timestamp 1696677024
transform 1 0 1548 0 -1 705
box -2 -3 26 103
use AND2X2  AND2X2_10
timestamp 1696677024
transform -1 0 1604 0 -1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_30
timestamp 1696677024
transform -1 0 1628 0 -1 705
box -2 -3 26 103
use NAND3X1  NAND3X1_18
timestamp 1696677024
transform -1 0 1660 0 -1 705
box -2 -3 34 103
use INVX2  INVX2_11
timestamp 1696677024
transform 1 0 1660 0 -1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_24
timestamp 1696677024
transform 1 0 1676 0 -1 705
box -2 -3 26 103
use INVX2  INVX2_10
timestamp 1696677024
transform 1 0 1700 0 -1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_51
timestamp 1696677024
transform -1 0 1740 0 -1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_40
timestamp 1696677024
transform -1 0 1772 0 -1 705
box -2 -3 34 103
use NOR2X1  NOR2X1_52
timestamp 1696677024
transform -1 0 1796 0 -1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_100
timestamp 1696677024
transform 1 0 1796 0 -1 705
box -2 -3 98 103
use BUFX2  BUFX2_23
timestamp 1696677024
transform 1 0 1892 0 -1 705
box -2 -3 26 103
use BUFX2  BUFX2_30
timestamp 1696677024
transform 1 0 1916 0 -1 705
box -2 -3 26 103
use FILL  FILL_7_1
timestamp 1696677024
transform -1 0 1948 0 -1 705
box -2 -3 10 103
use FILL  FILL_7_2
timestamp 1696677024
transform -1 0 1956 0 -1 705
box -2 -3 10 103
use CLKBUF1  CLKBUF1_18
timestamp 1696677024
transform 1 0 4 0 1 705
box -2 -3 74 103
use NOR2X1  NOR2X1_19
timestamp 1696677024
transform -1 0 100 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_48
timestamp 1696677024
transform -1 0 196 0 1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_38
timestamp 1696677024
transform 1 0 196 0 1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_25
timestamp 1696677024
transform 1 0 292 0 1 705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_94
timestamp 1696677024
transform -1 0 412 0 1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_40
timestamp 1696677024
transform 1 0 412 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_5
timestamp 1696677024
transform 1 0 436 0 1 705
box -2 -3 26 103
use FILL  FILL_7_0_0
timestamp 1696677024
transform -1 0 468 0 1 705
box -2 -3 10 103
use FILL  FILL_7_0_1
timestamp 1696677024
transform -1 0 476 0 1 705
box -2 -3 10 103
use NOR2X1  NOR2X1_32
timestamp 1696677024
transform -1 0 500 0 1 705
box -2 -3 26 103
use INVX1  INVX1_10
timestamp 1696677024
transform -1 0 516 0 1 705
box -2 -3 18 103
use NAND2X1  NAND2X1_10
timestamp 1696677024
transform -1 0 540 0 1 705
box -2 -3 26 103
use OAI21X1  OAI21X1_14
timestamp 1696677024
transform -1 0 572 0 1 705
box -2 -3 34 103
use OR2X2  OR2X2_2
timestamp 1696677024
transform 1 0 572 0 1 705
box -2 -3 34 103
use AOI21X1  AOI21X1_10
timestamp 1696677024
transform 1 0 604 0 1 705
box -2 -3 34 103
use NAND3X1  NAND3X1_4
timestamp 1696677024
transform -1 0 668 0 1 705
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_95
timestamp 1696677024
transform -1 0 764 0 1 705
box -2 -3 98 103
use AOI21X1  AOI21X1_11
timestamp 1696677024
transform 1 0 764 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_13
timestamp 1696677024
transform 1 0 796 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_15
timestamp 1696677024
transform -1 0 860 0 1 705
box -2 -3 34 103
use OAI21X1  OAI21X1_17
timestamp 1696677024
transform -1 0 892 0 1 705
box -2 -3 34 103
use BUFX4  BUFX4_14
timestamp 1696677024
transform -1 0 924 0 1 705
box -2 -3 34 103
use MUX2X1  MUX2X1_28
timestamp 1696677024
transform -1 0 972 0 1 705
box -2 -3 50 103
use FILL  FILL_7_1_0
timestamp 1696677024
transform 1 0 972 0 1 705
box -2 -3 10 103
use FILL  FILL_7_1_1
timestamp 1696677024
transform 1 0 980 0 1 705
box -2 -3 10 103
use BUFX4  BUFX4_6
timestamp 1696677024
transform 1 0 988 0 1 705
box -2 -3 34 103
use INVX8  INVX8_1
timestamp 1696677024
transform -1 0 1060 0 1 705
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_147
timestamp 1696677024
transform 1 0 1060 0 1 705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_133
timestamp 1696677024
transform 1 0 1156 0 1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_81
timestamp 1696677024
transform -1 0 1276 0 1 705
box -2 -3 26 103
use CLKBUF1  CLKBUF1_10
timestamp 1696677024
transform 1 0 1276 0 1 705
box -2 -3 74 103
use INVX8  INVX8_2
timestamp 1696677024
transform -1 0 1388 0 1 705
box -2 -3 42 103
use DFFPOSX1  DFFPOSX1_108
timestamp 1696677024
transform 1 0 1388 0 1 705
box -2 -3 98 103
use FILL  FILL_7_2_0
timestamp 1696677024
transform 1 0 1484 0 1 705
box -2 -3 10 103
use FILL  FILL_7_2_1
timestamp 1696677024
transform 1 0 1492 0 1 705
box -2 -3 10 103
use BUFX2  BUFX2_46
timestamp 1696677024
transform 1 0 1500 0 1 705
box -2 -3 26 103
use INVX1  INVX1_59
timestamp 1696677024
transform 1 0 1524 0 1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_98
timestamp 1696677024
transform 1 0 1540 0 1 705
box -2 -3 98 103
use NOR2X1  NOR2X1_53
timestamp 1696677024
transform -1 0 1660 0 1 705
box -2 -3 26 103
use NAND2X1  NAND2X1_25
timestamp 1696677024
transform 1 0 1660 0 1 705
box -2 -3 26 103
use INVX1  INVX1_21
timestamp 1696677024
transform 1 0 1684 0 1 705
box -2 -3 18 103
use OAI21X1  OAI21X1_41
timestamp 1696677024
transform -1 0 1732 0 1 705
box -2 -3 34 103
use INVX1  INVX1_20
timestamp 1696677024
transform 1 0 1732 0 1 705
box -2 -3 18 103
use NOR2X1  NOR2X1_50
timestamp 1696677024
transform -1 0 1772 0 1 705
box -2 -3 26 103
use AOI21X1  AOI21X1_26
timestamp 1696677024
transform -1 0 1804 0 1 705
box -2 -3 34 103
use NAND2X1  NAND2X1_26
timestamp 1696677024
transform -1 0 1828 0 1 705
box -2 -3 26 103
use INVX1  INVX1_22
timestamp 1696677024
transform -1 0 1844 0 1 705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_104
timestamp 1696677024
transform 1 0 1844 0 1 705
box -2 -3 98 103
use FILL  FILL_8_1
timestamp 1696677024
transform 1 0 1940 0 1 705
box -2 -3 10 103
use FILL  FILL_8_2
timestamp 1696677024
transform 1 0 1948 0 1 705
box -2 -3 10 103
use NAND2X1  NAND2X1_45
timestamp 1696677024
transform 1 0 4 0 -1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_8
timestamp 1696677024
transform -1 0 76 0 -1 905
box -2 -3 50 103
use MUX2X1  MUX2X1_6
timestamp 1696677024
transform 1 0 76 0 -1 905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_92
timestamp 1696677024
transform -1 0 220 0 -1 905
box -2 -3 98 103
use BUFX4  BUFX4_9
timestamp 1696677024
transform -1 0 252 0 -1 905
box -2 -3 34 103
use BUFX4  BUFX4_8
timestamp 1696677024
transform 1 0 252 0 -1 905
box -2 -3 34 103
use INVX2  INVX2_2
timestamp 1696677024
transform 1 0 284 0 -1 905
box -2 -3 18 103
use NOR2X1  NOR2X1_39
timestamp 1696677024
transform -1 0 324 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_17
timestamp 1696677024
transform 1 0 324 0 -1 905
box -2 -3 26 103
use INVX1  INVX1_7
timestamp 1696677024
transform 1 0 348 0 -1 905
box -2 -3 18 103
use NAND2X1  NAND2X1_7
timestamp 1696677024
transform 1 0 364 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_33
timestamp 1696677024
transform 1 0 388 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_12
timestamp 1696677024
transform -1 0 444 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_31
timestamp 1696677024
transform 1 0 444 0 -1 905
box -2 -3 26 103
use FILL  FILL_8_0_0
timestamp 1696677024
transform 1 0 468 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_0_1
timestamp 1696677024
transform 1 0 476 0 -1 905
box -2 -3 10 103
use XOR2X1  XOR2X1_2
timestamp 1696677024
transform 1 0 484 0 -1 905
box -2 -3 58 103
use OAI21X1  OAI21X1_48
timestamp 1696677024
transform -1 0 572 0 -1 905
box -2 -3 34 103
use INVX1  INVX1_37
timestamp 1696677024
transform -1 0 588 0 -1 905
box -2 -3 18 103
use NAND3X1  NAND3X1_3
timestamp 1696677024
transform 1 0 588 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_56
timestamp 1696677024
transform -1 0 716 0 -1 905
box -2 -3 98 103
use NAND2X1  NAND2X1_37
timestamp 1696677024
transform -1 0 740 0 -1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_40
timestamp 1696677024
transform -1 0 836 0 -1 905
box -2 -3 98 103
use BUFX4  BUFX4_5
timestamp 1696677024
transform -1 0 868 0 -1 905
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_55
timestamp 1696677024
transform -1 0 964 0 -1 905
box -2 -3 98 103
use FILL  FILL_8_1_0
timestamp 1696677024
transform -1 0 972 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_1_1
timestamp 1696677024
transform -1 0 980 0 -1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_134
timestamp 1696677024
transform -1 0 1076 0 -1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_150
timestamp 1696677024
transform -1 0 1172 0 -1 905
box -2 -3 98 103
use NOR2X1  NOR2X1_83
timestamp 1696677024
transform 1 0 1172 0 -1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_40
timestamp 1696677024
transform -1 0 1220 0 -1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_31
timestamp 1696677024
transform 1 0 1220 0 -1 905
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_59
timestamp 1696677024
transform -1 0 1364 0 -1 905
box -2 -3 98 103
use NOR2X1  NOR2X1_14
timestamp 1696677024
transform 1 0 1364 0 -1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_3
timestamp 1696677024
transform -1 0 1436 0 -1 905
box -2 -3 50 103
use FILL  FILL_8_2_0
timestamp 1696677024
transform -1 0 1444 0 -1 905
box -2 -3 10 103
use FILL  FILL_8_2_1
timestamp 1696677024
transform -1 0 1452 0 -1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_43
timestamp 1696677024
transform -1 0 1548 0 -1 905
box -2 -3 98 103
use BUFX2  BUFX2_51
timestamp 1696677024
transform 1 0 1548 0 -1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_66
timestamp 1696677024
transform 1 0 1572 0 -1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_55
timestamp 1696677024
transform -1 0 1628 0 -1 905
box -2 -3 26 103
use NAND3X1  NAND3X1_17
timestamp 1696677024
transform -1 0 1660 0 -1 905
box -2 -3 34 103
use NAND3X1  NAND3X1_16
timestamp 1696677024
transform 1 0 1660 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_49
timestamp 1696677024
transform 1 0 1692 0 -1 905
box -2 -3 26 103
use INVX2  INVX2_12
timestamp 1696677024
transform 1 0 1716 0 -1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_42
timestamp 1696677024
transform 1 0 1732 0 -1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_55
timestamp 1696677024
transform 1 0 1764 0 -1 905
box -2 -3 26 103
use NOR2X1  NOR2X1_54
timestamp 1696677024
transform -1 0 1812 0 -1 905
box -2 -3 26 103
use XNOR2X1  XNOR2X1_6
timestamp 1696677024
transform -1 0 1868 0 -1 905
box -2 -3 58 103
use BUFX2  BUFX2_35
timestamp 1696677024
transform -1 0 1892 0 -1 905
box -2 -3 26 103
use BUFX2  BUFX2_40
timestamp 1696677024
transform 1 0 1892 0 -1 905
box -2 -3 26 103
use BUFX2  BUFX2_12
timestamp 1696677024
transform 1 0 1916 0 -1 905
box -2 -3 26 103
use FILL  FILL_9_1
timestamp 1696677024
transform -1 0 1948 0 -1 905
box -2 -3 10 103
use FILL  FILL_9_2
timestamp 1696677024
transform -1 0 1956 0 -1 905
box -2 -3 10 103
use BUFX2  BUFX2_1
timestamp 1696677024
transform -1 0 28 0 1 905
box -2 -3 26 103
use OAI21X1  OAI21X1_59
timestamp 1696677024
transform -1 0 60 0 1 905
box -2 -3 34 103
use INVX1  INVX1_50
timestamp 1696677024
transform -1 0 76 0 1 905
box -2 -3 18 103
use XOR2X1  XOR2X1_5
timestamp 1696677024
transform 1 0 76 0 1 905
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_76
timestamp 1696677024
transform -1 0 228 0 1 905
box -2 -3 98 103
use NOR3X1  NOR3X1_11
timestamp 1696677024
transform -1 0 292 0 1 905
box -2 -3 66 103
use AOI21X1  AOI21X1_25
timestamp 1696677024
transform -1 0 324 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_38
timestamp 1696677024
transform 1 0 324 0 1 905
box -2 -3 34 103
use OAI21X1  OAI21X1_11
timestamp 1696677024
transform 1 0 356 0 1 905
box -2 -3 34 103
use NOR2X1  NOR2X1_85
timestamp 1696677024
transform -1 0 412 0 1 905
box -2 -3 26 103
use NAND2X1  NAND2X1_32
timestamp 1696677024
transform -1 0 436 0 1 905
box -2 -3 26 103
use AOI21X1  AOI21X1_9
timestamp 1696677024
transform -1 0 468 0 1 905
box -2 -3 34 103
use FILL  FILL_9_0_0
timestamp 1696677024
transform -1 0 476 0 1 905
box -2 -3 10 103
use FILL  FILL_9_0_1
timestamp 1696677024
transform -1 0 484 0 1 905
box -2 -3 10 103
use XNOR2X1  XNOR2X1_1
timestamp 1696677024
transform -1 0 540 0 1 905
box -2 -3 58 103
use NAND2X1  NAND2X1_36
timestamp 1696677024
transform -1 0 564 0 1 905
box -2 -3 26 103
use NOR3X1  NOR3X1_9
timestamp 1696677024
transform 1 0 564 0 1 905
box -2 -3 66 103
use XOR2X1  XOR2X1_1
timestamp 1696677024
transform -1 0 684 0 1 905
box -2 -3 58 103
use INVX1  INVX1_38
timestamp 1696677024
transform 1 0 684 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_49
timestamp 1696677024
transform 1 0 700 0 1 905
box -2 -3 34 103
use MUX2X1  MUX2X1_16
timestamp 1696677024
transform 1 0 732 0 1 905
box -2 -3 50 103
use NOR2X1  NOR2X1_27
timestamp 1696677024
transform -1 0 804 0 1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_15
timestamp 1696677024
transform 1 0 804 0 1 905
box -2 -3 50 103
use NOR2X1  NOR2X1_26
timestamp 1696677024
transform -1 0 876 0 1 905
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_39
timestamp 1696677024
transform -1 0 972 0 1 905
box -2 -3 98 103
use FILL  FILL_9_1_0
timestamp 1696677024
transform 1 0 972 0 1 905
box -2 -3 10 103
use FILL  FILL_9_1_1
timestamp 1696677024
transform 1 0 980 0 1 905
box -2 -3 10 103
use CLKBUF1  CLKBUF1_5
timestamp 1696677024
transform 1 0 988 0 1 905
box -2 -3 74 103
use NOR2X1  NOR2X1_84
timestamp 1696677024
transform 1 0 1060 0 1 905
box -2 -3 26 103
use MUX2X1  MUX2X1_32
timestamp 1696677024
transform 1 0 1084 0 1 905
box -2 -3 50 103
use OAI21X1  OAI21X1_54
timestamp 1696677024
transform -1 0 1164 0 1 905
box -2 -3 34 103
use NAND2X1  NAND2X1_41
timestamp 1696677024
transform -1 0 1188 0 1 905
box -2 -3 26 103
use INVX1  INVX1_44
timestamp 1696677024
transform -1 0 1204 0 1 905
box -2 -3 18 103
use OAI21X1  OAI21X1_53
timestamp 1696677024
transform -1 0 1236 0 1 905
box -2 -3 34 103
use INVX1  INVX1_43
timestamp 1696677024
transform -1 0 1252 0 1 905
box -2 -3 18 103
use XOR2X1  XOR2X1_3
timestamp 1696677024
transform -1 0 1308 0 1 905
box -2 -3 58 103
use NOR3X1  NOR3X1_10
timestamp 1696677024
transform 1 0 1308 0 1 905
box -2 -3 66 103
use XOR2X1  XOR2X1_4
timestamp 1696677024
transform 1 0 1372 0 1 905
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_72
timestamp 1696677024
transform -1 0 1524 0 1 905
box -2 -3 98 103
use FILL  FILL_9_2_0
timestamp 1696677024
transform -1 0 1532 0 1 905
box -2 -3 10 103
use FILL  FILL_9_2_1
timestamp 1696677024
transform -1 0 1540 0 1 905
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_88
timestamp 1696677024
transform -1 0 1636 0 1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_102
timestamp 1696677024
transform 1 0 1636 0 1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_99
timestamp 1696677024
transform -1 0 1828 0 1 905
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_103
timestamp 1696677024
transform 1 0 1828 0 1 905
box -2 -3 98 103
use BUFX2  BUFX2_33
timestamp 1696677024
transform 1 0 1924 0 1 905
box -2 -3 26 103
use FILL  FILL_10_1
timestamp 1696677024
transform 1 0 1948 0 1 905
box -2 -3 10 103
use NAND2X1  NAND2X1_43
timestamp 1696677024
transform 1 0 4 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_57
timestamp 1696677024
transform -1 0 60 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_48
timestamp 1696677024
transform -1 0 76 0 -1 1105
box -2 -3 18 103
use AND2X2  AND2X2_16
timestamp 1696677024
transform 1 0 76 0 -1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_95
timestamp 1696677024
transform 1 0 108 0 -1 1105
box -2 -3 26 103
use OAI22X1  OAI22X1_3
timestamp 1696677024
transform -1 0 172 0 -1 1105
box -2 -3 42 103
use NAND2X1  NAND2X1_42
timestamp 1696677024
transform 1 0 172 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_56
timestamp 1696677024
transform -1 0 228 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_47
timestamp 1696677024
transform -1 0 244 0 -1 1105
box -2 -3 18 103
use XOR2X1  XOR2X1_6
timestamp 1696677024
transform 1 0 244 0 -1 1105
box -2 -3 58 103
use NAND2X1  NAND2X1_44
timestamp 1696677024
transform 1 0 300 0 -1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_58
timestamp 1696677024
transform -1 0 356 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_49
timestamp 1696677024
transform -1 0 372 0 -1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_19
timestamp 1696677024
transform 1 0 372 0 -1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_15
timestamp 1696677024
transform 1 0 396 0 -1 1105
box -2 -3 34 103
use FILL  FILL_10_0_0
timestamp 1696677024
transform 1 0 428 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_0_1
timestamp 1696677024
transform 1 0 436 0 -1 1105
box -2 -3 10 103
use NOR3X1  NOR3X1_4
timestamp 1696677024
transform 1 0 444 0 -1 1105
box -2 -3 66 103
use BUFX4  BUFX4_12
timestamp 1696677024
transform -1 0 540 0 -1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_14
timestamp 1696677024
transform 1 0 540 0 -1 1105
box -2 -3 50 103
use NAND2X1  NAND2X1_35
timestamp 1696677024
transform 1 0 588 0 -1 1105
box -2 -3 26 103
use OAI22X1  OAI22X1_1
timestamp 1696677024
transform 1 0 612 0 -1 1105
box -2 -3 42 103
use NOR2X1  NOR2X1_87
timestamp 1696677024
transform 1 0 652 0 -1 1105
box -2 -3 26 103
use AND2X2  AND2X2_12
timestamp 1696677024
transform 1 0 676 0 -1 1105
box -2 -3 34 103
use OAI21X1  OAI21X1_47
timestamp 1696677024
transform -1 0 740 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_36
timestamp 1696677024
transform -1 0 756 0 -1 1105
box -2 -3 18 103
use CLKBUF1  CLKBUF1_3
timestamp 1696677024
transform -1 0 828 0 -1 1105
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_120
timestamp 1696677024
transform -1 0 924 0 -1 1105
box -2 -3 98 103
use FILL  FILL_10_1_0
timestamp 1696677024
transform -1 0 932 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_1_1
timestamp 1696677024
transform -1 0 940 0 -1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_136
timestamp 1696677024
transform -1 0 1036 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_148
timestamp 1696677024
transform -1 0 1132 0 -1 1105
box -2 -3 98 103
use NOR2X1  NOR2X1_82
timestamp 1696677024
transform 1 0 1132 0 -1 1105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_1
timestamp 1696677024
transform -1 0 1228 0 -1 1105
box -2 -3 74 103
use MUX2X1  MUX2X1_29
timestamp 1696677024
transform 1 0 1228 0 -1 1105
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_71
timestamp 1696677024
transform 1 0 1276 0 -1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_87
timestamp 1696677024
transform 1 0 1372 0 -1 1105
box -2 -3 98 103
use NAND2X1  NAND2X1_38
timestamp 1696677024
transform 1 0 1468 0 -1 1105
box -2 -3 26 103
use FILL  FILL_10_2_0
timestamp 1696677024
transform -1 0 1500 0 -1 1105
box -2 -3 10 103
use FILL  FILL_10_2_1
timestamp 1696677024
transform -1 0 1508 0 -1 1105
box -2 -3 10 103
use OAI21X1  OAI21X1_51
timestamp 1696677024
transform -1 0 1540 0 -1 1105
box -2 -3 34 103
use INVX1  INVX1_41
timestamp 1696677024
transform -1 0 1556 0 -1 1105
box -2 -3 18 103
use NOR2X1  NOR2X1_91
timestamp 1696677024
transform 1 0 1556 0 -1 1105
box -2 -3 26 103
use OAI22X1  OAI22X1_2
timestamp 1696677024
transform -1 0 1620 0 -1 1105
box -2 -3 42 103
use NOR2X1  NOR2X1_90
timestamp 1696677024
transform 1 0 1620 0 -1 1105
box -2 -3 26 103
use AND2X2  AND2X2_13
timestamp 1696677024
transform -1 0 1676 0 -1 1105
box -2 -3 34 103
use MUX2X1  MUX2X1_1
timestamp 1696677024
transform 1 0 1676 0 -1 1105
box -2 -3 50 103
use NOR2X1  NOR2X1_12
timestamp 1696677024
transform -1 0 1748 0 -1 1105
box -2 -3 26 103
use CLKBUF1  CLKBUF1_2
timestamp 1696677024
transform 1 0 1748 0 -1 1105
box -2 -3 74 103
use MUX2X1  MUX2X1_38
timestamp 1696677024
transform -1 0 1868 0 -1 1105
box -2 -3 50 103
use MUX2X1  MUX2X1_40
timestamp 1696677024
transform 1 0 1868 0 -1 1105
box -2 -3 50 103
use OR2X2  OR2X2_7
timestamp 1696677024
transform 1 0 1916 0 -1 1105
box -2 -3 34 103
use FILL  FILL_11_1
timestamp 1696677024
transform -1 0 1956 0 -1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_90
timestamp 1696677024
transform -1 0 100 0 1 1105
box -2 -3 98 103
use NOR2X1  NOR2X1_94
timestamp 1696677024
transform 1 0 100 0 1 1105
box -2 -3 26 103
use AND2X2  AND2X2_15
timestamp 1696677024
transform 1 0 124 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_68
timestamp 1696677024
transform 1 0 156 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_84
timestamp 1696677024
transform -1 0 348 0 1 1105
box -2 -3 98 103
use OAI21X1  OAI21X1_32
timestamp 1696677024
transform 1 0 348 0 1 1105
box -2 -3 34 103
use AOI21X1  AOI21X1_21
timestamp 1696677024
transform -1 0 412 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_41
timestamp 1696677024
transform 1 0 412 0 1 1105
box -2 -3 26 103
use NAND3X1  NAND3X1_12
timestamp 1696677024
transform -1 0 468 0 1 1105
box -2 -3 34 103
use FILL  FILL_11_0_0
timestamp 1696677024
transform -1 0 476 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_0_1
timestamp 1696677024
transform -1 0 484 0 1 1105
box -2 -3 10 103
use NAND3X1  NAND3X1_9
timestamp 1696677024
transform -1 0 516 0 1 1105
box -2 -3 34 103
use NAND3X1  NAND3X1_10
timestamp 1696677024
transform -1 0 548 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_14
timestamp 1696677024
transform -1 0 564 0 1 1105
box -2 -3 18 103
use NAND2X1  NAND2X1_16
timestamp 1696677024
transform -1 0 588 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_31
timestamp 1696677024
transform -1 0 620 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_13
timestamp 1696677024
transform -1 0 636 0 1 1105
box -2 -3 18 103
use AND2X2  AND2X2_11
timestamp 1696677024
transform -1 0 668 0 1 1105
box -2 -3 34 103
use NOR2X1  NOR2X1_86
timestamp 1696677024
transform 1 0 668 0 1 1105
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_66
timestamp 1696677024
transform -1 0 788 0 1 1105
box -2 -3 98 103
use INVX1  INVX1_35
timestamp 1696677024
transform -1 0 804 0 1 1105
box -2 -3 18 103
use OAI21X1  OAI21X1_46
timestamp 1696677024
transform 1 0 804 0 1 1105
box -2 -3 34 103
use NAND2X1  NAND2X1_34
timestamp 1696677024
transform -1 0 860 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_26
timestamp 1696677024
transform 1 0 860 0 1 1105
box -2 -3 50 103
use NOR2X1  NOR2X1_78
timestamp 1696677024
transform -1 0 932 0 1 1105
box -2 -3 26 103
use FILL  FILL_11_1_0
timestamp 1696677024
transform -1 0 940 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_1_1
timestamp 1696677024
transform -1 0 948 0 1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_132
timestamp 1696677024
transform -1 0 1044 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_42
timestamp 1696677024
transform 1 0 1044 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_58
timestamp 1696677024
transform -1 0 1236 0 1 1105
box -2 -3 98 103
use NOR2X1  NOR2X1_13
timestamp 1696677024
transform 1 0 1236 0 1 1105
box -2 -3 26 103
use MUX2X1  MUX2X1_2
timestamp 1696677024
transform -1 0 1308 0 1 1105
box -2 -3 50 103
use NAND2X1  NAND2X1_4
timestamp 1696677024
transform -1 0 1332 0 1 1105
box -2 -3 26 103
use NOR2X1  NOR2X1_28
timestamp 1696677024
transform 1 0 1332 0 1 1105
box -2 -3 26 103
use NAND2X1  NAND2X1_39
timestamp 1696677024
transform 1 0 1356 0 1 1105
box -2 -3 26 103
use OAI21X1  OAI21X1_52
timestamp 1696677024
transform -1 0 1412 0 1 1105
box -2 -3 34 103
use INVX1  INVX1_42
timestamp 1696677024
transform -1 0 1428 0 1 1105
box -2 -3 18 103
use INVX1  INVX1_8
timestamp 1696677024
transform -1 0 1444 0 1 1105
box -2 -3 18 103
use FILL  FILL_11_2_0
timestamp 1696677024
transform -1 0 1452 0 1 1105
box -2 -3 10 103
use FILL  FILL_11_2_1
timestamp 1696677024
transform -1 0 1460 0 1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_41
timestamp 1696677024
transform -1 0 1556 0 1 1105
box -2 -3 98 103
use AND2X2  AND2X2_14
timestamp 1696677024
transform 1 0 1556 0 1 1105
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_57
timestamp 1696677024
transform -1 0 1684 0 1 1105
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_86
timestamp 1696677024
transform -1 0 1780 0 1 1105
box -2 -3 98 103
use MUX2X1  MUX2X1_39
timestamp 1696677024
transform -1 0 1828 0 1 1105
box -2 -3 50 103
use OAI21X1  OAI21X1_55
timestamp 1696677024
transform -1 0 1860 0 1 1105
box -2 -3 34 103
use BUFX2  BUFX2_11
timestamp 1696677024
transform 1 0 1860 0 1 1105
box -2 -3 26 103
use AOI21X1  AOI21X1_34
timestamp 1696677024
transform 1 0 1884 0 1 1105
box -2 -3 34 103
use BUFX2  BUFX2_37
timestamp 1696677024
transform 1 0 1916 0 1 1105
box -2 -3 26 103
use FILL  FILL_12_1
timestamp 1696677024
transform 1 0 1940 0 1 1105
box -2 -3 10 103
use FILL  FILL_12_2
timestamp 1696677024
transform 1 0 1948 0 1 1105
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_74
timestamp 1696677024
transform -1 0 100 0 -1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_130
timestamp 1696677024
transform -1 0 196 0 -1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_146
timestamp 1696677024
transform 1 0 196 0 -1 1305
box -2 -3 98 103
use INVX2  INVX2_6
timestamp 1696677024
transform 1 0 292 0 -1 1305
box -2 -3 18 103
use NAND2X1  NAND2X1_18
timestamp 1696677024
transform 1 0 308 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_16
timestamp 1696677024
transform 1 0 332 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_37
timestamp 1696677024
transform -1 0 380 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_37
timestamp 1696677024
transform 1 0 380 0 -1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_8
timestamp 1696677024
transform -1 0 436 0 -1 1305
box -2 -3 34 103
use INVX1  INVX1_15
timestamp 1696677024
transform 1 0 436 0 -1 1305
box -2 -3 18 103
use FILL  FILL_12_0_0
timestamp 1696677024
transform -1 0 460 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_0_1
timestamp 1696677024
transform -1 0 468 0 -1 1305
box -2 -3 10 103
use OAI21X1  OAI21X1_34
timestamp 1696677024
transform -1 0 500 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_38
timestamp 1696677024
transform -1 0 524 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_17
timestamp 1696677024
transform 1 0 524 0 -1 1305
box -2 -3 18 103
use NAND3X1  NAND3X1_14
timestamp 1696677024
transform 1 0 540 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_43
timestamp 1696677024
transform 1 0 572 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_15
timestamp 1696677024
transform -1 0 620 0 -1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_14
timestamp 1696677024
transform -1 0 644 0 -1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_6
timestamp 1696677024
transform -1 0 676 0 -1 1305
box -2 -3 34 103
use NOR2X1  NOR2X1_36
timestamp 1696677024
transform -1 0 700 0 -1 1305
box -2 -3 26 103
use NOR3X1  NOR3X1_3
timestamp 1696677024
transform 1 0 700 0 -1 1305
box -2 -3 66 103
use NOR2X1  NOR2X1_42
timestamp 1696677024
transform 1 0 764 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_26
timestamp 1696677024
transform 1 0 788 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_13
timestamp 1696677024
transform -1 0 844 0 -1 1305
box -2 -3 26 103
use INVX4  INVX4_1
timestamp 1696677024
transform 1 0 844 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_35
timestamp 1696677024
transform 1 0 868 0 -1 1305
box -2 -3 26 103
use INVX1  INVX1_12
timestamp 1696677024
transform -1 0 908 0 -1 1305
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_82
timestamp 1696677024
transform -1 0 1004 0 -1 1305
box -2 -3 98 103
use FILL  FILL_12_1_0
timestamp 1696677024
transform -1 0 1012 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_1_1
timestamp 1696677024
transform -1 0 1020 0 -1 1305
box -2 -3 10 103
use CLKBUF1  CLKBUF1_16
timestamp 1696677024
transform -1 0 1092 0 -1 1305
box -2 -3 74 103
use BUFX4  BUFX4_10
timestamp 1696677024
transform -1 0 1124 0 -1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_30
timestamp 1696677024
transform 1 0 1124 0 -1 1305
box -2 -3 50 103
use INVX1  INVX1_40
timestamp 1696677024
transform 1 0 1172 0 -1 1305
box -2 -3 18 103
use BUFX4  BUFX4_1
timestamp 1696677024
transform -1 0 1220 0 -1 1305
box -2 -3 34 103
use CLKBUF1  CLKBUF1_11
timestamp 1696677024
transform 1 0 1220 0 -1 1305
box -2 -3 74 103
use BUFX4  BUFX4_4
timestamp 1696677024
transform 1 0 1292 0 -1 1305
box -2 -3 34 103
use BUFX4  BUFX4_13
timestamp 1696677024
transform 1 0 1324 0 -1 1305
box -2 -3 34 103
use INVX2  INVX2_3
timestamp 1696677024
transform -1 0 1372 0 -1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_22
timestamp 1696677024
transform 1 0 1372 0 -1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_15
timestamp 1696677024
transform -1 0 1436 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_6
timestamp 1696677024
transform 1 0 1436 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_30
timestamp 1696677024
transform 1 0 1460 0 -1 1305
box -2 -3 26 103
use FILL  FILL_12_2_0
timestamp 1696677024
transform -1 0 1492 0 -1 1305
box -2 -3 10 103
use FILL  FILL_12_2_1
timestamp 1696677024
transform -1 0 1500 0 -1 1305
box -2 -3 10 103
use NOR2X1  NOR2X1_29
timestamp 1696677024
transform -1 0 1524 0 -1 1305
box -2 -3 26 103
use AOI21X1  AOI21X1_14
timestamp 1696677024
transform 1 0 1524 0 -1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_2
timestamp 1696677024
transform -1 0 1588 0 -1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_3
timestamp 1696677024
transform -1 0 1612 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_34
timestamp 1696677024
transform -1 0 1636 0 -1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_20
timestamp 1696677024
transform -1 0 1668 0 -1 1305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_2
timestamp 1696677024
transform -1 0 1724 0 -1 1305
box -2 -3 58 103
use DFFPOSX1  DFFPOSX1_70
timestamp 1696677024
transform -1 0 1820 0 -1 1305
box -2 -3 98 103
use MUX2X1  MUX2X1_37
timestamp 1696677024
transform -1 0 1868 0 -1 1305
box -2 -3 50 103
use INVX1  INVX1_52
timestamp 1696677024
transform 1 0 1868 0 -1 1305
box -2 -3 18 103
use NOR2X1  NOR2X1_92
timestamp 1696677024
transform 1 0 1884 0 -1 1305
box -2 -3 26 103
use BUFX2  BUFX2_10
timestamp 1696677024
transform 1 0 1908 0 -1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_93
timestamp 1696677024
transform 1 0 1932 0 -1 1305
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_63
timestamp 1696677024
transform -1 0 100 0 1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_47
timestamp 1696677024
transform 1 0 100 0 1 1305
box -2 -3 98 103
use NOR2X1  NOR2X1_18
timestamp 1696677024
transform 1 0 196 0 1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_7
timestamp 1696677024
transform 1 0 220 0 1 1305
box -2 -3 50 103
use BUFX2  BUFX2_45
timestamp 1696677024
transform 1 0 268 0 1 1305
box -2 -3 26 103
use NOR2X1  NOR2X1_72
timestamp 1696677024
transform -1 0 316 0 1 1305
box -2 -3 26 103
use MUX2X1  MUX2X1_20
timestamp 1696677024
transform -1 0 364 0 1 1305
box -2 -3 50 103
use OAI21X1  OAI21X1_35
timestamp 1696677024
transform -1 0 396 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_23
timestamp 1696677024
transform -1 0 428 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_13
timestamp 1696677024
transform 1 0 428 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_0_0
timestamp 1696677024
transform -1 0 468 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_0_1
timestamp 1696677024
transform -1 0 476 0 1 1305
box -2 -3 10 103
use XNOR2X1  XNOR2X1_4
timestamp 1696677024
transform -1 0 532 0 1 1305
box -2 -3 58 103
use BUFX4  BUFX4_11
timestamp 1696677024
transform -1 0 564 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_28
timestamp 1696677024
transform 1 0 564 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_29
timestamp 1696677024
transform -1 0 628 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_5
timestamp 1696677024
transform 1 0 628 0 1 1305
box -2 -3 34 103
use NAND3X1  NAND3X1_11
timestamp 1696677024
transform 1 0 660 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_9
timestamp 1696677024
transform 1 0 692 0 1 1305
box -2 -3 26 103
use NAND3X1  NAND3X1_7
timestamp 1696677024
transform 1 0 716 0 1 1305
box -2 -3 34 103
use XNOR2X1  XNOR2X1_3
timestamp 1696677024
transform 1 0 748 0 1 1305
box -2 -3 58 103
use MUX2X1  MUX2X1_27
timestamp 1696677024
transform 1 0 804 0 1 1305
box -2 -3 50 103
use AOI21X1  AOI21X1_19
timestamp 1696677024
transform 1 0 852 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_27
timestamp 1696677024
transform -1 0 916 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_34
timestamp 1696677024
transform -1 0 964 0 1 1305
box -2 -3 50 103
use FILL  FILL_13_1_0
timestamp 1696677024
transform -1 0 972 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_1_1
timestamp 1696677024
transform -1 0 980 0 1 1305
box -2 -3 10 103
use BUFX4  BUFX4_3
timestamp 1696677024
transform -1 0 1012 0 1 1305
box -2 -3 34 103
use MUX2X1  MUX2X1_45
timestamp 1696677024
transform 1 0 1012 0 1 1305
box -2 -3 50 103
use MUX2X1  MUX2X1_46
timestamp 1696677024
transform -1 0 1108 0 1 1305
box -2 -3 50 103
use INVX1  INVX1_58
timestamp 1696677024
transform 1 0 1108 0 1 1305
box -2 -3 18 103
use MUX2X1  MUX2X1_47
timestamp 1696677024
transform -1 0 1172 0 1 1305
box -2 -3 50 103
use MUX2X1  MUX2X1_48
timestamp 1696677024
transform 1 0 1172 0 1 1305
box -2 -3 50 103
use MUX2X1  MUX2X1_25
timestamp 1696677024
transform -1 0 1268 0 1 1305
box -2 -3 50 103
use MUX2X1  MUX2X1_4
timestamp 1696677024
transform 1 0 1268 0 1 1305
box -2 -3 50 103
use AOI21X1  AOI21X1_16
timestamp 1696677024
transform -1 0 1348 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_23
timestamp 1696677024
transform 1 0 1348 0 1 1305
box -2 -3 34 103
use OR2X2  OR2X2_3
timestamp 1696677024
transform -1 0 1412 0 1 1305
box -2 -3 34 103
use NAND2X1  NAND2X1_12
timestamp 1696677024
transform -1 0 1436 0 1 1305
box -2 -3 26 103
use NAND2X1  NAND2X1_11
timestamp 1696677024
transform 1 0 1436 0 1 1305
box -2 -3 26 103
use OAI21X1  OAI21X1_21
timestamp 1696677024
transform -1 0 1492 0 1 1305
box -2 -3 34 103
use FILL  FILL_13_2_0
timestamp 1696677024
transform 1 0 1492 0 1 1305
box -2 -3 10 103
use FILL  FILL_13_2_1
timestamp 1696677024
transform 1 0 1500 0 1 1305
box -2 -3 10 103
use INVX1  INVX1_11
timestamp 1696677024
transform 1 0 1508 0 1 1305
box -2 -3 18 103
use OAI21X1  OAI21X1_19
timestamp 1696677024
transform 1 0 1524 0 1 1305
box -2 -3 34 103
use INVX2  INVX2_4
timestamp 1696677024
transform 1 0 1556 0 1 1305
box -2 -3 18 103
use AOI21X1  AOI21X1_17
timestamp 1696677024
transform 1 0 1572 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_24
timestamp 1696677024
transform 1 0 1604 0 1 1305
box -2 -3 34 103
use OAI21X1  OAI21X1_18
timestamp 1696677024
transform -1 0 1668 0 1 1305
box -2 -3 34 103
use AOI21X1  AOI21X1_13
timestamp 1696677024
transform -1 0 1700 0 1 1305
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_69
timestamp 1696677024
transform 1 0 1700 0 1 1305
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_85
timestamp 1696677024
transform -1 0 1892 0 1 1305
box -2 -3 98 103
use BUFX2  BUFX2_9
timestamp 1696677024
transform 1 0 1892 0 1 1305
box -2 -3 26 103
use BUFX2  BUFX2_13
timestamp 1696677024
transform 1 0 1916 0 1 1305
box -2 -3 26 103
use FILL  FILL_14_1
timestamp 1696677024
transform 1 0 1940 0 1 1305
box -2 -3 10 103
use FILL  FILL_14_2
timestamp 1696677024
transform 1 0 1948 0 1 1305
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_45
timestamp 1696677024
transform -1 0 100 0 -1 1505
box -2 -3 98 103
use NOR2X1  NOR2X1_16
timestamp 1696677024
transform 1 0 100 0 -1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_5
timestamp 1696677024
transform 1 0 124 0 -1 1505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_73
timestamp 1696677024
transform -1 0 268 0 -1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_89
timestamp 1696677024
transform -1 0 364 0 -1 1505
box -2 -3 98 103
use OAI21X1  OAI21X1_36
timestamp 1696677024
transform -1 0 396 0 -1 1505
box -2 -3 34 103
use AOI21X1  AOI21X1_24
timestamp 1696677024
transform -1 0 428 0 -1 1505
box -2 -3 34 103
use INVX2  INVX2_7
timestamp 1696677024
transform 1 0 428 0 -1 1505
box -2 -3 18 103
use FILL  FILL_14_0_0
timestamp 1696677024
transform -1 0 452 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_0_1
timestamp 1696677024
transform -1 0 460 0 -1 1505
box -2 -3 10 103
use XNOR2X1  XNOR2X1_5
timestamp 1696677024
transform -1 0 516 0 -1 1505
box -2 -3 58 103
use AOI21X1  AOI21X1_22
timestamp 1696677024
transform 1 0 516 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_33
timestamp 1696677024
transform -1 0 580 0 -1 1505
box -2 -3 34 103
use INVX2  INVX2_5
timestamp 1696677024
transform 1 0 580 0 -1 1505
box -2 -3 18 103
use AOI21X1  AOI21X1_20
timestamp 1696677024
transform 1 0 596 0 -1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_18
timestamp 1696677024
transform 1 0 628 0 -1 1505
box -2 -3 50 103
use BUFX4  BUFX4_2
timestamp 1696677024
transform -1 0 708 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_30
timestamp 1696677024
transform -1 0 740 0 -1 1505
box -2 -3 34 103
use DFFPOSX1  DFFPOSX1_121
timestamp 1696677024
transform -1 0 836 0 -1 1505
box -2 -3 98 103
use NOR2X1  NOR2X1_79
timestamp 1696677024
transform 1 0 836 0 -1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_18
timestamp 1696677024
transform 1 0 860 0 -1 1505
box -2 -3 34 103
use OAI21X1  OAI21X1_25
timestamp 1696677024
transform -1 0 924 0 -1 1505
box -2 -3 34 103
use MUX2X1  MUX2X1_35
timestamp 1696677024
transform -1 0 972 0 -1 1505
box -2 -3 50 103
use FILL  FILL_14_1_0
timestamp 1696677024
transform 1 0 972 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_1_1
timestamp 1696677024
transform 1 0 980 0 -1 1505
box -2 -3 10 103
use MUX2X1  MUX2X1_33
timestamp 1696677024
transform 1 0 988 0 -1 1505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_135
timestamp 1696677024
transform -1 0 1132 0 -1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_119
timestamp 1696677024
transform -1 0 1228 0 -1 1505
box -2 -3 98 103
use NOR2X1  NOR2X1_77
timestamp 1696677024
transform -1 0 1252 0 -1 1505
box -2 -3 26 103
use CLKBUF1  CLKBUF1_17
timestamp 1696677024
transform -1 0 1324 0 -1 1505
box -2 -3 74 103
use DFFPOSX1  DFFPOSX1_60
timestamp 1696677024
transform -1 0 1420 0 -1 1505
box -2 -3 98 103
use CLKBUF1  CLKBUF1_15
timestamp 1696677024
transform 1 0 1420 0 -1 1505
box -2 -3 74 103
use FILL  FILL_14_2_0
timestamp 1696677024
transform 1 0 1492 0 -1 1505
box -2 -3 10 103
use FILL  FILL_14_2_1
timestamp 1696677024
transform 1 0 1500 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_143
timestamp 1696677024
transform 1 0 1508 0 -1 1505
box -2 -3 98 103
use NAND2X1  NAND2X1_20
timestamp 1696677024
transform 1 0 1604 0 -1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_23
timestamp 1696677024
transform 1 0 1628 0 -1 1505
box -2 -3 50 103
use NOR2X1  NOR2X1_44
timestamp 1696677024
transform -1 0 1700 0 -1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_75
timestamp 1696677024
transform -1 0 1724 0 -1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_125
timestamp 1696677024
transform 1 0 1724 0 -1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_141
timestamp 1696677024
transform 1 0 1820 0 -1 1505
box -2 -3 98 103
use BUFX2  BUFX2_42
timestamp 1696677024
transform 1 0 1916 0 -1 1505
box -2 -3 26 103
use FILL  FILL_15_1
timestamp 1696677024
transform -1 0 1948 0 -1 1505
box -2 -3 10 103
use FILL  FILL_15_2
timestamp 1696677024
transform -1 0 1956 0 -1 1505
box -2 -3 10 103
use DFFPOSX1  DFFPOSX1_61
timestamp 1696677024
transform -1 0 100 0 1 1505
box -2 -3 98 103
use MUX2X1  MUX2X1_42
timestamp 1696677024
transform -1 0 148 0 1 1505
box -2 -3 50 103
use BUFX2  BUFX2_20
timestamp 1696677024
transform -1 0 28 0 -1 1705
box -2 -3 26 103
use BUFX2  BUFX2_21
timestamp 1696677024
transform -1 0 52 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_97
timestamp 1696677024
transform -1 0 76 0 -1 1705
box -2 -3 26 103
use INVX1  INVX1_51
timestamp 1696677024
transform -1 0 92 0 -1 1705
box -2 -3 18 103
use OAI21X1  OAI21X1_60
timestamp 1696677024
transform 1 0 92 0 -1 1705
box -2 -3 34 103
use MUX2X1  MUX2X1_43
timestamp 1696677024
transform -1 0 196 0 1 1505
box -2 -3 50 103
use MUX2X1  MUX2X1_41
timestamp 1696677024
transform -1 0 244 0 1 1505
box -2 -3 50 103
use AOI21X1  AOI21X1_35
timestamp 1696677024
transform -1 0 156 0 -1 1705
box -2 -3 34 103
use BUFX2  BUFX2_19
timestamp 1696677024
transform 1 0 156 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_96
timestamp 1696677024
transform -1 0 204 0 -1 1705
box -2 -3 26 103
use BUFX2  BUFX2_18
timestamp 1696677024
transform 1 0 204 0 -1 1705
box -2 -3 26 103
use MUX2X1  MUX2X1_44
timestamp 1696677024
transform -1 0 292 0 1 1505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_91
timestamp 1696677024
transform -1 0 388 0 1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_145
timestamp 1696677024
transform -1 0 324 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_75
timestamp 1696677024
transform 1 0 388 0 1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_129
timestamp 1696677024
transform -1 0 420 0 -1 1705
box -2 -3 98 103
use FILL  FILL_15_0_0
timestamp 1696677024
transform -1 0 492 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_0_1
timestamp 1696677024
transform -1 0 500 0 1 1505
box -2 -3 10 103
use INVX1  INVX1_46
timestamp 1696677024
transform -1 0 516 0 1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_71
timestamp 1696677024
transform 1 0 420 0 -1 1705
box -2 -3 26 103
use FILL  FILL_16_0_0
timestamp 1696677024
transform 1 0 444 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_0_1
timestamp 1696677024
transform 1 0 452 0 -1 1705
box -2 -3 10 103
use MUX2X1  MUX2X1_19
timestamp 1696677024
transform 1 0 460 0 -1 1705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_144
timestamp 1696677024
transform -1 0 604 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_83
timestamp 1696677024
transform -1 0 612 0 1 1505
box -2 -3 98 103
use NOR2X1  NOR2X1_70
timestamp 1696677024
transform -1 0 628 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_67
timestamp 1696677024
transform -1 0 708 0 1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_65
timestamp 1696677024
transform -1 0 804 0 1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_128
timestamp 1696677024
transform -1 0 724 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_81
timestamp 1696677024
transform -1 0 900 0 1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_137
timestamp 1696677024
transform -1 0 820 0 -1 1705
box -2 -3 98 103
use MUX2X1  MUX2X1_36
timestamp 1696677024
transform -1 0 948 0 1 1505
box -2 -3 50 103
use BUFX2  BUFX2_4
timestamp 1696677024
transform -1 0 844 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_89
timestamp 1696677024
transform 1 0 844 0 -1 1705
box -2 -3 26 103
use BUFX2  BUFX2_5
timestamp 1696677024
transform -1 0 892 0 -1 1705
box -2 -3 26 103
use INVX1  INVX1_39
timestamp 1696677024
transform -1 0 908 0 -1 1705
box -2 -3 18 103
use DFFPOSX1  DFFPOSX1_53
timestamp 1696677024
transform -1 0 1004 0 -1 1705
box -2 -3 98 103
use AOI21X1  AOI21X1_33
timestamp 1696677024
transform 1 0 948 0 1 1505
box -2 -3 34 103
use FILL  FILL_15_1_0
timestamp 1696677024
transform 1 0 980 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_1_1
timestamp 1696677024
transform 1 0 988 0 1 1505
box -2 -3 10 103
use OAI21X1  OAI21X1_50
timestamp 1696677024
transform 1 0 996 0 1 1505
box -2 -3 34 103
use FILL  FILL_16_1_0
timestamp 1696677024
transform 1 0 1004 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_1_1
timestamp 1696677024
transform 1 0 1012 0 -1 1705
box -2 -3 10 103
use NOR2X1  NOR2X1_88
timestamp 1696677024
transform -1 0 1052 0 1 1505
box -2 -3 26 103
use BUFX2  BUFX2_2
timestamp 1696677024
transform 1 0 1052 0 1 1505
box -2 -3 26 103
use BUFX2  BUFX2_3
timestamp 1696677024
transform 1 0 1076 0 1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_13
timestamp 1696677024
transform 1 0 1100 0 1 1505
box -2 -3 50 103
use NOR2X1  NOR2X1_24
timestamp 1696677024
transform 1 0 1020 0 -1 1705
box -2 -3 26 103
use BUFX2  BUFX2_8
timestamp 1696677024
transform 1 0 1044 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_37
timestamp 1696677024
transform -1 0 1164 0 -1 1705
box -2 -3 98 103
use BUFX2  BUFX2_26
timestamp 1696677024
transform -1 0 1172 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_100
timestamp 1696677024
transform 1 0 1172 0 1 1505
box -2 -3 26 103
use AOI21X1  AOI21X1_36
timestamp 1696677024
transform -1 0 1228 0 1 1505
box -2 -3 34 103
use BUFX2  BUFX2_27
timestamp 1696677024
transform -1 0 1188 0 -1 1705
box -2 -3 26 103
use BUFX2  BUFX2_29
timestamp 1696677024
transform 1 0 1188 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_142
timestamp 1696677024
transform -1 0 1308 0 -1 1705
box -2 -3 98 103
use OAI21X1  OAI21X1_65
timestamp 1696677024
transform -1 0 1260 0 1 1505
box -2 -3 34 103
use INVX1  INVX1_57
timestamp 1696677024
transform 1 0 1260 0 1 1505
box -2 -3 18 103
use NOR2X1  NOR2X1_101
timestamp 1696677024
transform 1 0 1276 0 1 1505
box -2 -3 26 103
use BUFX2  BUFX2_28
timestamp 1696677024
transform 1 0 1300 0 1 1505
box -2 -3 26 103
use BUFX2  BUFX2_6
timestamp 1696677024
transform -1 0 1332 0 -1 1705
box -2 -3 26 103
use NOR2X1  NOR2X1_15
timestamp 1696677024
transform -1 0 1348 0 1 1505
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_44
timestamp 1696677024
transform -1 0 1444 0 1 1505
box -2 -3 98 103
use BUFX2  BUFX2_15
timestamp 1696677024
transform 1 0 1332 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_126
timestamp 1696677024
transform 1 0 1356 0 -1 1705
box -2 -3 98 103
use MUX2X1  MUX2X1_17
timestamp 1696677024
transform -1 0 1492 0 1 1505
box -2 -3 50 103
use FILL  FILL_15_2_0
timestamp 1696677024
transform -1 0 1500 0 1 1505
box -2 -3 10 103
use FILL  FILL_15_2_1
timestamp 1696677024
transform -1 0 1508 0 1 1505
box -2 -3 10 103
use NOR2X1  NOR2X1_69
timestamp 1696677024
transform -1 0 1532 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_76
timestamp 1696677024
transform 1 0 1452 0 -1 1705
box -2 -3 26 103
use FILL  FILL_16_2_0
timestamp 1696677024
transform 1 0 1476 0 -1 1705
box -2 -3 10 103
use FILL  FILL_16_2_1
timestamp 1696677024
transform 1 0 1484 0 -1 1705
box -2 -3 10 103
use MUX2X1  MUX2X1_24
timestamp 1696677024
transform 1 0 1492 0 -1 1705
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_127
timestamp 1696677024
transform 1 0 1532 0 1 1505
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_123
timestamp 1696677024
transform -1 0 1636 0 -1 1705
box -2 -3 98 103
use AND2X2  AND2X2_3
timestamp 1696677024
transform -1 0 1660 0 1 1505
box -2 -3 34 103
use NOR2X1  NOR2X1_73
timestamp 1696677024
transform 1 0 1660 0 1 1505
box -2 -3 26 103
use MUX2X1  MUX2X1_21
timestamp 1696677024
transform -1 0 1732 0 1 1505
box -2 -3 50 103
use DFFPOSX1  DFFPOSX1_139
timestamp 1696677024
transform 1 0 1636 0 -1 1705
box -2 -3 98 103
use MUX2X1  MUX2X1_22
timestamp 1696677024
transform 1 0 1732 0 1 1505
box -2 -3 50 103
use BUFX2  BUFX2_43
timestamp 1696677024
transform -1 0 1804 0 1 1505
box -2 -3 26 103
use NOR2X1  NOR2X1_74
timestamp 1696677024
transform -1 0 1828 0 1 1505
box -2 -3 26 103
use BUFX2  BUFX2_22
timestamp 1696677024
transform 1 0 1732 0 -1 1705
box -2 -3 26 103
use DFFPOSX1  DFFPOSX1_140
timestamp 1696677024
transform -1 0 1852 0 -1 1705
box -2 -3 98 103
use DFFPOSX1  DFFPOSX1_124
timestamp 1696677024
transform 1 0 1828 0 1 1505
box -2 -3 98 103
use BUFX2  BUFX2_16
timestamp 1696677024
transform -1 0 1876 0 -1 1705
box -2 -3 26 103
use BUFX2  BUFX2_14
timestamp 1696677024
transform 1 0 1876 0 -1 1705
box -2 -3 26 103
use BUFX2  BUFX2_7
timestamp 1696677024
transform 1 0 1900 0 -1 1705
box -2 -3 26 103
use BUFX2  BUFX2_31
timestamp 1696677024
transform 1 0 1924 0 1 1505
box -2 -3 26 103
use FILL  FILL_16_1
timestamp 1696677024
transform 1 0 1948 0 1 1505
box -2 -3 10 103
use INVX1  INVX1_26
timestamp 1696677024
transform 1 0 1924 0 -1 1705
box -2 -3 18 103
use FILL  FILL_17_1
timestamp 1696677024
transform -1 0 1948 0 -1 1705
box -2 -3 10 103
use FILL  FILL_17_2
timestamp 1696677024
transform -1 0 1956 0 -1 1705
box -2 -3 10 103
<< labels >>
flabel metal6 s 456 -30 472 -22 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal6 s 968 -30 984 -22 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 654 -22 658 -18 7 FreeSans 24 270 0 0 clock
port 2 nsew
flabel metal2 s 1702 1728 1706 1732 3 FreeSans 24 90 0 0 key[0]
port 3 nsew
flabel metal2 s 1758 1728 1762 1732 3 FreeSans 24 90 0 0 key[1]
port 4 nsew
flabel metal2 s 1678 1728 1682 1732 3 FreeSans 24 90 0 0 key[2]
port 5 nsew
flabel metal2 s 1510 1728 1514 1732 3 FreeSans 24 90 0 0 key[3]
port 6 nsew
flabel metal3 s -26 738 -22 742 7 FreeSans 24 0 0 0 reset
port 7 nsew
flabel metal3 s -26 248 -22 252 7 FreeSans 24 0 0 0 time_button
port 8 nsew
flabel metal2 s 766 -22 770 -18 7 FreeSans 24 270 0 0 alarm_button
port 9 nsew
flabel metal3 s 1982 848 1986 852 3 FreeSans 24 0 0 0 fastwatch
port 10 nsew
flabel metal2 s 214 1728 218 1732 3 FreeSans 24 90 0 0 ms_hour[0]
port 11 nsew
flabel metal2 s 166 1728 170 1732 3 FreeSans 24 90 0 0 ms_hour[1]
port 12 nsew
flabel metal3 s -26 1668 -22 1672 7 FreeSans 24 90 0 0 ms_hour[2]
port 13 nsew
flabel metal3 s -26 1648 -22 1652 7 FreeSans 24 90 0 0 ms_hour[3]
port 14 nsew
flabel metal2 s 1742 1728 1746 1732 3 FreeSans 24 90 0 0 ms_hour[4]
port 15 nsew
flabel metal3 s 1982 648 1986 652 3 FreeSans 24 0 0 0 ms_hour[5]
port 16 nsew
flabel metal3 s -26 648 -22 652 7 FreeSans 24 0 0 0 ms_hour[6]
port 17 nsew
flabel metal3 s -26 448 -22 452 7 FreeSans 24 0 0 0 ms_hour[7]
port 18 nsew
flabel metal2 s 1062 1728 1066 1732 3 FreeSans 24 90 0 0 ls_hour[0]
port 19 nsew
flabel metal2 s 1094 1728 1098 1732 3 FreeSans 24 90 0 0 ls_hour[1]
port 20 nsew
flabel metal2 s 830 1728 834 1732 3 FreeSans 24 90 0 0 ls_hour[2]
port 21 nsew
flabel metal2 s 878 1728 882 1732 3 FreeSans 24 90 0 0 ls_hour[3]
port 22 nsew
flabel metal2 s 1310 1728 1314 1732 3 FreeSans 24 90 0 0 ls_hour[4]
port 23 nsew
flabel metal2 s 1910 1728 1914 1732 3 FreeSans 24 90 0 0 ls_hour[5]
port 24 nsew
flabel metal2 s 1078 1728 1082 1732 3 FreeSans 24 90 0 0 ls_hour[6]
port 25 nsew
flabel metal3 s 1982 1368 1986 1372 3 FreeSans 24 0 0 0 ls_hour[7]
port 26 nsew
flabel metal2 s 1158 1728 1162 1732 3 FreeSans 24 90 0 0 ms_minute[0]
port 27 nsew
flabel metal2 s 1174 1728 1178 1732 3 FreeSans 24 90 0 0 ms_minute[1]
port 28 nsew
flabel metal2 s 1326 1728 1330 1732 3 FreeSans 24 90 0 0 ms_minute[2]
port 29 nsew
flabel metal2 s 1198 1728 1202 1732 3 FreeSans 24 90 0 0 ms_minute[3]
port 30 nsew
flabel metal3 s 1982 668 1986 672 3 FreeSans 24 0 0 0 ms_minute[4]
port 31 nsew
flabel metal3 s 1982 1548 1986 1552 3 FreeSans 24 0 0 0 ms_minute[5]
port 32 nsew
flabel metal2 s 574 -22 578 -18 7 FreeSans 24 270 0 0 ms_minute[6]
port 33 nsew
flabel metal3 s 1982 948 1986 952 3 FreeSans 24 0 0 0 ms_minute[7]
port 34 nsew
flabel metal3 s 1982 1248 1986 1252 3 FreeSans 24 0 0 0 ls_minute[0]
port 35 nsew
flabel metal3 s 1982 1148 1986 1152 3 FreeSans 24 0 0 0 ls_minute[1]
port 36 nsew
flabel metal3 s 1982 868 1986 872 3 FreeSans 24 0 0 0 ls_minute[2]
port 37 nsew
flabel metal3 s 1982 1348 1986 1352 3 FreeSans 24 0 0 0 ls_minute[3]
port 38 nsew
flabel metal2 s 1886 1728 1890 1732 3 FreeSans 24 90 0 0 ls_minute[4]
port 39 nsew
flabel metal2 s 1342 1728 1346 1732 3 FreeSans 24 90 0 0 ls_minute[5]
port 40 nsew
flabel metal2 s 1862 1728 1866 1732 3 FreeSans 24 90 0 0 ls_minute[6]
port 41 nsew
flabel metal3 s -26 148 -22 152 7 FreeSans 24 0 0 0 ls_minute[7]
port 42 nsew
flabel metal3 s -26 948 -22 952 7 FreeSans 24 0 0 0 alarm_sound
port 43 nsew
<< end >>
